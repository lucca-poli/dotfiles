Vim�UnDo� F�B��8�E~�P�F�\�8j2v�Lܑ�\?g�  Y                                   f�    _�                             ����                                                                                                                                                                                                                                                                                                                                                             f�     �              5��                                                5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f�     �               5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f�    �               5��                                                  5�_�                     :        ����                                                                                                                                                                                                                                                                                                                                                  V        f�     �   9   ;        5��    9                      �                     5��