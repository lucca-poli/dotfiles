Vim�UnDo� O��f��`��J%��V�}s�vq���q���}��   P   .    signal count : integer;  -- Input stimulus                            f��    _�                     	       ����                                                                                                                                                                                                                                                                                                                                      	          V       f�l     �         M    �   	   
   M    �      	          C            clk : in bit;                            -- Clock input   A            rst : in bit;                          -- Reset input   F            count : out integer       -- 6-bit count output (64 steps)5��                          �       �               �                          �               �       5�_�                    	       ����                                                                                                                                                                                                                                                                                                                            	                           f�p    �   	      P              done: out bit;   O        count : out unsigned(5 downto 0)       -- 6-bit count output (64 steps)�      
   P      C        clk, rst: in bit;                            -- Clock input5��                         �                      �    	                     �                      �    
                                          5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         P      .    signal count : integer;  -- Input stimulus5��                        (                    �                         *                     �                         )                     �                        (                    �                         *                     �                         )                     �                        (                    �                        (                    �                         *                     �                         )                     �                        (                    �                        (                    �                        (                    �                        (                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f��    �         P      ;    signal count : unsigned(7 downto 0);  -- Input stimulus5��                        1                    5�_�                    >       ����                                                                                                                                                                                                                                                                                                                                                v       f��    �   >   ?   P    �   >   ?   P              wait for CLOCK_PERIOD;5��    >                      �                     5�_�                    ?       ����                                                                                                                                                                                                                                                                                                                                                v       f��     �   ?   @   Q    �   ?   @   Q              wait for CLOCK_PERIOD;5��    ?                      �                     5�_�                    @       ����                                                                                                                                                                                                                                                                                                                                                v       f��     �   @   A   R    �   @   A   R              wait for CLOCK_PERIOD;5��    @                      �                     5�_�      	              A       ����                                                                                                                                                                                                                                                                                                                                                v       f��     �   A   B   S    �   A   B   S              wait for CLOCK_PERIOD;5��    A                      �                     5�_�      
           	   B       ����                                                                                                                                                                                                                                                                                                                                                v       f��     �   B   C   T    �   B   C   T              wait for CLOCK_PERIOD;5��    B                                           5�_�   	              
   C       ����                                                                                                                                                                                                                                                                                                                                                v       f��     �   C   D   U    �   C   D   U              wait for CLOCK_PERIOD;5��    C                      "                     5�_�   
                  D       ����                                                                                                                                                                                                                                                                                                                                                v       f��    �   D   E   V    �   D   E   V              wait for CLOCK_PERIOD;5��    D                      A                     5��