Vim�UnDo� &�r�ƅ�g��,
U���WZ�K_)�*�   5           wait;   2         !      !   !       f��    _�                             ����                                                                                                                                                                                                                                                                                                                                                             f�i     �                   �               5��                    @                       �      5�_�                    	        ����                                                                                                                                                                                                                                                                                                                            	                      V        f�     �         =    �   	   
   =    �      	                      clk, rst : in bit;   /            msgi : in bit_vector(511 downto 0);   0            haso : out bit_vector(255 downto 0);               done : out bit5��                          �       �               �                          �               1       5�_�                    	       ����                                                                                                                                                                                                                                                                                                                            	          
                 f�     �   	      ?              clk_out: out bit�      
   ?              clk_in: in bit;5��                         �                      �    	                     �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                            	          
                 f�     �         ?      entity multisteps_tb is end;5��              
          *       
              5�_�                           ����                                                                                                                                                                                                                                                                                                                            	          
                 f�     �         ?      +architecture Behavioral of multisteps_tb is5��                        Z                     �                         \                      �                         [                      �                        Z                     �                        Z                     �                        Z                     5�_�                       %    ����                                                                                                                                                                                                                                                                                                                            	          
                 f�     �                -    signal rst : bit := '0';  -- Reset signal5��                          c      .               5�_�                            ����                                                                                                                                                                                                                                                                                                                            	          
                 f�     �                Q    signal msgi : bit_vector(511 downto 0) := (others => '0');  -- Input stimulus5��                          w      R               5�_�      	                      ����                                                                                                                                                                                                                                                                                                                            	          
                 f�     �                >    signal haso : bit_vector(255 downto 0);  -- Input stimulus5��                          w      ?               5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                            	          
                 f�     �         <          signal done: bit;5��                        �                    5�_�   	              
   "   	    ����                                                                                                                                                                                                                                                                                                                            	          
                 f��     �   !   #   <          dut: multisteps5��    !   	       
          �      
              �    !                     �                     �    !   
                  �                     �    !   	                 �                    �    !                     �                     �    !                     �                     �    !                     �                     �    !                     �                     �    !                     �                     �    !   
                  �                     �    !   	                 �                    �    !                     �                     �    !                     �                     �    !                     �                     �    !                     �                     �    !                     �                     �    !                     �                     �    !                     �                     �    !                     �                     �    !                     �                     �    !   
                  �                     �    !   	                 �                    �    !   	                 �                    �    !   	                 �                    5�_�   
                        ����                                                                                                                                                                                                                                                                                                                            	          
                 f��     �         <          component multisteps5��              
          w       
              �                        w                     �                        w                     �                        w                     �                        w                     �                        w                     �                                               5�_�                    "       ����                                                                                                                                                                                                                                                                                                                            	          
                 f��     �   !   #   <          dut: slow_clk_tb5��    !                     �                     5�_�                    "       ����                                                                                                                                                                                                                                                                                                                            	          
                 f��     �   !   #   <          dut: slow_clk_t5��    !                     �                     5�_�                    "       ����                                                                                                                                                                                                                                                                                                                            	          
                 f��     �   !   #   <          dut: slow_clk_5��    !                     �                     5�_�                    $       ����                                                                                                                                                                                                                                                                                                                            	          
                 f��     �   #   $                      clk => clk,5��    #                      �                     5�_�                    $       ����                                                                                                                                                                                                                                                                                                                            	          
                 f��     �   #   $                      rst => rst,5��    #                      �                     5�_�                    $       ����                                                                                                                                                                                                                                                                                                                            	          
                 f��     �   #   $                      msgi => msgi,5��    #                      �                     5�_�                    $       ����                                                                                                                                                                                                                                                                                                                            	          
                 f��     �   #   %   9                  haso => haso,5��    #                     �                     �    #                     �                    5�_�                    %       ����                                                                                                                                                                                                                                                                                                                            	          
                 f��     �   $   &   9                  done => done5��    $                    �                    �    $                     �                     �    $                     �                     �    $                    �                    �    $                    �                    �    $                    �                    5�_�                    .       ����                                                                                                                                                                                                                                                                                                                            	          
                 f�     �   -   .                  if done = '1' then5��    -                      p                     5�_�                    .       ����                                                                                                                                                                                                                                                                                                                            	          
                 f�     �   -   .                      assert false report5��    -                      p                      5�_�                    .       ����                                                                                                                                                                                                                                                                                                                            	          
                 f�     �   -   .          (            "haso = " & to_hstring(haso)5��    -                      p      )               5�_�                    .       ����                                                                                                                                                                                                                                                                                                                            	          
                 f�     �   -   .                      severity note;5��    -                      p                     5�_�                    .       ����                                                                                                                                                                                                                                                                                                                            	          
                 f�     �   -   /   5              end if;5��    -                    x                    �    -   
                  z                     �    -   	                  y                     �    -                    x                    �    -                    x                    �    -                 
   x             
       �    -                    �                    �    -                    �                    �    -                     �                     �    -                    �                    �    -                     �                     �    -                     �                     5�_�                    .       ����                                                                                                                                                                                                                                                                                                                            	          
                 f�*     �   -   /   5              wait for 15��    -                     �                     5�_�                    .       ����                                                                                                                                                                                                                                                                                                                            	          
                 f�3    �   -   /   5              wait for 1ms;5��    -                     �                     5�_�                    0   !    ����                                                                                                                                                                                                                                                                                                                            	          
                 f�     �   /   1   5      ;        assert false report "EOT multisteps" severity note;5��    /   !       
          �      
              5�_�                    ,   !    ����                                                                                                                                                                                                                                                                                                                            	          
                 f�    �   +   -   5      ;        assert false report "BOT multisteps" severity note;5��    +   !       
          T      
              �    +   !                 T                    5�_�                   2       ����                                                                                                                                                                                                                                                                                                                            	          
                 f��     �   1   3   5              wait for 1s;5��    1                     �                     5�_�                     2       ����                                                                                                                                                                                                                                                                                                                            	          
                 f��     �   1   3   5              wait for 1 s;5��    1                     �                     5�_�      !               2       ����                                                                                                                                                                                                                                                                                                                            	          
                 f��     �   1   3   5              wait for 1 ms;5��    1                     �                     5�_�                   !   2       ����                                                                                                                                                                                                                                                                                                                            	          
                 f��    �   1   3   5              wait for 10 ms;5��    1                     �                     5�_�                    2       ����                                                                                                                                                                                                                                                                                                                            	          
                 f��    �   1   3        5��    1                      �                     5��