Vim�UnDo� �\��@"���},)�ɧ@��s�����&s$��     ,    signal contagem: bit_vector(3 downto 0);   �                           f)FG    _�                            ����                                                                                                                                                                                                                                                                                                                                                             f)D�     �   �   �          ?      -- clockRecepcao: divisorclock4 port map(clock, '0', CR);�   �   �          >      clockTransmissao: divisorclock port map(clock, '0', CT);�   Y   [                component divisorclock is�   S   U          #      -- component divisorclock4 is�                '    architecture arc of divisorclock is�   	                 end divisorclock;�                  entity divisorclock is5��                        X                     �    	                    �                     �                        	                    �    S                    �	                    �    Y                    .
                    �    �                                        �    �                    N                    5�_�                    �        ����                                                                                                                                                                                                                                                                                                                                                             f)D�     �   �   �        ?      clockTransmissao: clock_divider port map(clock, '0', CT);5��    �                    �                    5�_�                    1        ����                                                                                                                                                                                                                                                                                                                                                             f)E     �  q  s          �    REGISTRADORC: registrador_entrada_serial generic map(TAMANHO_REG => (WIDTH + 1)) port map(shift_sig, serial_data, registrador_out);�  8  :          ,    component registrador_entrada_serial is �  6  8          4    architecture serial_in_arch of entrada_serial is�  4  6              end entrada_serial ;�  (  *          entity entrada_serial is�   �   �          >architecture registrador_arch of registrador_entrada_serial is�   �   �          %entity registrador_entrada_serial is �   �   �          f      entrada_serialC: entrada_serial port map(CR, reset, '1', serial_in, done_SI, parity_SI, byteIn);�   0   2        !      component entrada_serial is5��    0                    h                    �    �                    �                    �    �                    �                    �    �                    ,%                    �    �   -                 0&                    �    (                   �+                    �    4                   -                    �    6  #                 ;-                    �    8                   �-                    �    q                   �9                    5�_�                   �        ����                                                                                                                                                                                                                                                                                                                                                             f)E-     �  q  s          �    REGISTRADORC: registrador_serial_input generic map(TAMANHO_REG => (WIDTH + 1)) port map(shift_sig, serial_data, registrador_out);�              (    end process ATUALIZACAO_REGISTRADOR;�   �   �        /    ATUALIZACAO_REGISTRADOR: process (shift) is5��    �                    �&                    �                       �'                    �    q                   �9                    5�_�      
            
        ����                                                                                                                                                                                                                                                                                                                                                             f)E<     �  s  u          k    CONTADOR10C: contador generic map(WIDTH => 4) port map(bit_sig, clr10_sig, enable_sig, contador10_out);�  r  t          f    CONTADOR4C: contador generic map(WIDTH => 3) port map(clock, clr4_sig, enable_sig, contador4_out);�  h  j          �    shift_sig <= not(contador4_out(2)) and contador4_out(1) and not contador4_out(0) when present_state = recebendo else '0'; --010 amostragem�  g  i          [    bit_sig <= contador4_out(2) and not(contador4_out(1)) and not(contador4_out(0)); --100 �  f  h          z    dado_sig_stop <= contador10_out(3) and contador10_out(2) and not(contador10_out(1)) and not(contador10_out(0)); --1100�  e  g          u    dado_sig <= contador10_out(3) and not(contador10_out(2)) and contador10_out(1) and not(contador10_out(0)); --1010�  U  W          2    signal contador10_out: bit_vector(3 downto 0);�  T  V          1    signal contador4_out: bit_vector(2 downto 0);�  C  E              component contador is�  !  #                  end contador64_arch;�              /    architecture contador64_arch of contador is�  	               entity contador is5��    	                   (                    �                       )                    �      #                 *)                    �    !                   �*                    �    C                   x.                    �    T                   ;1                    �    U                   l1                    �    e                   �5                    �    e  )                 �5                    �    e  ?                 �5                    �    e  X                 �5                    �    f                   *6                    �    f  *                 ?6                    �    f  C                 X6                    �    f  ]                 r6                    �    g                   �6                    �    g  '                 �6                    �    g  @                 �6                    �    h                   �6                    �    h  *                 7                    �    h  B                 '7                    �    r                   :                    �    r  V                 W:                    �    s                   w:                    �    s  Z                 �:                    5�_�         	       
   �        ����                                                                                                                                                                                                                                                                                                                                                             f)EP     �  q  s          �    REGISTERC: registrador_serial_input generic map(TAMANHO_REG => (WIDTH + 1)) port map(shift_sig, serial_data, registrador_out);�  ?  A          3        q: out bit_vector(TAMANHO_REG - 1 downto 0)�  :  <          !        TAMANHO_REG: natural := 9�   �            /            q_signal(TAMANHO_REG-1) <= data_in;�   �             Q            q_signal(TAMANHO_REG-2 downto 0) <= q_signal(TAMANHO_REG-1 downto 1);�   �   �          4signal q_signal: bit_vector(TAMANHO_REG-1 downto 0);�   �   �          1        q: out bit_vector(TAMANHO_REG-1 downto 0)�   �   �        1    TAMANHO_REG: natural := 9 -- 9 btis no total 5��    �                    N%                    �    �                    �%                    �    �                    V&                    �    �                    �&                    �    �   6                 '                    �    �                    D'                    �    :                   �-                    �    ?                   .                    �    q  4                 �9                    5�_�   
                s        ����                                                                                                                                                                                                                                                                                                                                                             f)E[     �  s  u          i    CONTADOR10C: counter generic map(WIDTH => 4) port map(bit_sig, clr10_sig, enable_sig, counter10_out);�  r  t        d    CONTADOR4C: counter generic map(WIDTH => 3) port map(clock, clr4_sig, enable_sig, counter4_out);5��    r                   �9                    �    s                   N:                    5�_�                   o        ����                                                                                                                                                                                                                                                                                                                                                             f)En     �  |  ~          8    estado_fim <= '1' when present_state = fim else '0';�  {  }          D    estado_recebendo <= '1' when present_state = recebendo else '0';�  z  |          N    estado_esperando_zero <= '1' when present_state = esperando_zero else '0';�  y  {          >    estado_inicio <= '1' when present_state = inicio else '0';�  [  ]              -- Máquina de estados�  V  X          p    signal estado_inicio, estado_esperando_zero, estado_recebendo, estado_fim, tick: bit; -- sinais para debugar�   n   p              --Maquina de estados5��    n                    9                    �    V                   �1                    �    V                   �1                    �    V  /                 �1                    �    V  @                 �1                    �    [                   3                    �    y                   �;                    �    z                   %<                    �    {                   s<                    �    |                   �<                    5�_�                    b        ����                                                                                                                                                                                                                                                                                                                                                             f)E|     �  y  {          =    state_inicio <= '1' when present_state = inicio else '0';�  l  n          5    clr4_sig <= '1' when present_state = inicio else �  k  m          :                 '1' when present_state = inicio else '0';�  ^  `          Q    next_state <= esperando_zero when present_state = inicio and start = '1' else�  \  ^          1    present_state <= inicio when reset = '1' else�  V  X          l    signal state_inicio, state_esperando_zero, state_recebendo, state_fim, tick: bit; -- sinais para debugar�  P  R          U    type state_type is (inicio, esperando_zero, recebendo, esperando_stop_bits, fim);�   q   s          m      next_state <= recebendo_dado when present_state = inicio and serial_in = '0' else -- recebe o start bit�   o   q          3      present_state <= inicio when reset = '1' else�   a   c        V      type state_type is (inicio, recebendo_dado, calculando, transmitindo_dado, fim);5��    a                                        �    o                    W                    �    q   8                 �                    �    P                   �/                    �    V                   �1                    �    \                   )3                    �    ^  6                 �3                    �    k  *                 8                    �    l  )                 P8                    �    y  
                 �;                    �    y  -                 <                    5�_�                   Q        ����                                                                                                                                                                                                                                                                                                                                                             f)E�     �  z  |          M    state_esperando_zero <= '1' when present_state = esperando_zero else '0';�  i  k          e    enable_sig <= '1' when present_state = recebendo or present_state = esperando_stop_bits else '0';�  b  d          K                  esperando_zero when present_state = fim and start = '1'; �  a  c          [                  fim when present_state = esperando_stop_bits and dado_sig_stop = '1' else�  `  b          \                  esperando_stop_bits when present_state = recebendo and dado_sig = '1' else�  _  a          W                  recebendo when present_state = esperando_zero and zero_sig = '1' else�  ^  `          Q    next_state <= esperando_zero when present_state = intial and start = '1' else�  V  X          l    signal state_intial, state_esperando_zero, state_recebendo, state_fim, tick: bit; -- sinais para debugar�  P  R        U    type state_type is (intial, esperando_zero, recebendo, esperando_stop_bits, fim);5��    P          	          �/      	              �    P  9       	          �/      	              �    V         	          �1      	              �    ^         	          �3      	              �    _  1       	          �3      	              �    `         	          14      	              �    a  +       	          �4      	              �    b         	          �4      	              �    i  H       	          �7      	              �    z  
       	          <      	              �    z  3       	          B<      	              5�_�                    b        ����                                                                                                                                                                                                                                                                                                                                                             f)E�     �  y  {          =    state_intial <= '1' when present_state = intial else '0';�  l  n          5    clr4_sig <= '1' when present_state = intial else �  k  m          :                 '1' when present_state = intial else '0';�  ^  `          O    next_state <= waiting_zero when present_state = intial and start = '1' else�  \  ^          1    present_state <= intial when reset = '1' else�  V  X          j    signal state_intial, state_waiting_zero, state_recebendo, state_fim, tick: bit; -- sinais para debugar�  P  R          Q    type state_type is (intial, waiting_zero, recebendo, waiting_stop_bits, fim);�   q   s          m      next_state <= recebendo_dado when present_state = intial and serial_in = '0' else -- recebe o start bit�   o   q          3      present_state <= intial when reset = '1' else�   a   c        V      type state_type is (intial, recebendo_dado, calculando, transmitindo_dado, fim);5��    a                                        �    o                    X                    �    q   8                 �                    �    P                   �/                    �    V                   �1                    �    \                   (3                    �    ^  4                 �3                    �    k  *                 8                    �    l  )                 F8                    �    y  
                 �;                    �    y  .                 <                    5�_�                    b        ����                                                                                                                                                                                                                                                                                                                                                             f)E�     �  {  }          C    state_recebendo <= '1' when present_state = recebendo else '0';�  i  k          c    enable_sig <= '1' when present_state = recebendo or present_state = waiting_stop_bits else '0';�  h  j          �    shift_sig <= not(counter4_out(2)) and counter4_out(1) and not counter4_out(0) when present_state = recebendo else '0'; --010 amostragem�  `  b          Z                  waiting_stop_bits when present_state = recebendo and dado_sig = '1' else�  _  a          U                  recebendo when present_state = waiting_zero and zero_sig = '1' else�  V  X          k    signal state_initial, state_waiting_zero, state_recebendo, state_fim, tick: bit; -- sinais para debugar�  P  R          R    type state_type is (initial, waiting_zero, recebendo, waiting_stop_bits, fim);�   v   x          X                    recebendo_dado when present_state = fim and serial_in = '0'; -- loop�   s   u          �                    recebendo_dado when present_state = calculando and serial_in = '0' else -- recebendo um dado no meio do caculo�   r   t          z                    calculando when present_state = recebendo_dado and done_SI = '1' else -- quando terminarmos de receber�   q   s          n      next_state <= recebendo_dado when present_state = initial and serial_in = '0' else -- recebe o start bit�   a   c        W      type state_type is (initial, recebendo_dado, calculando, transmitindo_dado, fim);5��    a   #       	       	   $      	       	       �    q          	       	   �      	       	       �    r   4       	       	   T      	       	       �    s          	       	   �      	       	       �    s   _       	       	   �      	       	       �    v          	       	   #      	       	       �    P  /       	       	   �/      	       	       �    V  4       	       	   �1      	       	       �    _         	       	   �3      	       	       �    `  9       	       	   _4      	       	       �    h  g       	       	   %7      	       	       �    i  +       	       	   u7      	       	       �    {  
       	       	   n<      	       	       �    {  0       	       	   �<      	       	       5�_�                   b        ����                                                                                                                                                                                                                                                                                                                                                             f)E�     �  |  ~          7    state_fim <= '1' when present_state = fim else '0';�  v  x          2    done <= '1' when present_state = fim else '0';�  u  w          L    parity_bit <= registrador_out((WIDTH + 1) - 1) when present_state = fim;�  j  l          2    clr10_sig <= '1' when present_state = fim else�  b  d          I                  waiting_zero when present_state = fim and start = '1'; �  a  c          Y                  fim when present_state = waiting_stop_bits and dado_sig_stop = '1' else�  V  X          k    signal state_initial, state_waiting_zero, state_receiving, state_fim, tick: bit; -- sinais para debugar�  P  R          R    type state_type is (initial, waiting_zero, receiving, waiting_stop_bits, fim);�   v   x          X                    receiving_dado when present_state = fim and serial_in = '0'; -- loop�   u   w          q                    fim when present_state = transmitindo_dado and done_SO = '1' else -- terminamos de trasnmitir�   a   c        W      type state_type is (initial, receiving_dado, calculando, transmitindo_dado, fim);5��    a   R                 S                    �    u                    �                    �    v   8                 K                    �    P  M                 0                    �    V  E                 �1                    �    a                   �4                    �    b  4                 5                    �    j  *                 �7                    �    u  H                 <;                    �    v  %                 h;                    �    |  
                 �<                    �    |  ,                 �<                    5�_�                   8       ����                                                                                                                                                                                                                                                                                                                                                             f)E�     �  7  9        .    -- Componentes ---------------------------5��    7                
   >-             
       5�_�                   &       ����                                                                                                                                                                                                                                                                                                                                                             f)E�     �  %  '        l----Top entidade -------------------------------------------------------------------------------------------5��    %                   )+                    5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f)E�     �   �   �        V-- entidades--------------------------------------------------------------------------5��    �          	          �$      	              5�_�                    �   
    ����                                                                                                                                                                                                                                                                                                                                                             f)F
     �   �   �              --sinais de auxilio--5��    �                      �                     5�_�                   O        ����                                                                                                                                                                                                                                                                                                                                                             f)F'     �  e  g          v    dado_sig_stop <= counter10_out(3) and counter10_out(2) and not(counter10_out(1)) and not(counter10_out(0)); --1100�  d  f          q    dado_sig <= counter10_out(3) and not(counter10_out(2)) and counter10_out(1) and not(counter10_out(0)); --1010�  b  d               -- Setting dados de controle�  `  b          [                  ended when present_state = waiting_stop_bits and dado_sig_stop = '1' else�  _  a          Z                  waiting_stop_bits when present_state = receiving and dado_sig = '1' else�  Q  S          s    signal serial_sig, shift_sig, zero_sig, enable_sig, bit_sig, dado_sig, dado_sig_stop, clr10_sig, clr4_sig: bit;�   �   �          K          serial_o <= data(to_integer(contagem_unsigned)-1); --saindo dados�   �   �          .    signal dado: bit_vector(WIDTH-1 downto 0);�   }             A      start_SO <= '1' when present_state = transmitindo_dado else�   {   }          A      reset_SO <= '0' when present_state = transmitindo_dado else�   v   x          Z                    receiving_dado when present_state = ended and serial_in = '0'; -- loop�   u   w          s                    ended when present_state = transmitindo_dado and done_SO = '1' else -- terminamos de trasnmitir�   t   v          ~                    transmitindo_dado when present_state = calculando and done_MS = '1' else -- quando terminarmos de calcular�   s   u          �                    receiving_dado when present_state = calculando and serial_in = '0' else -- receiving um dado no meio do caculo�   r   t          z                    calculando when present_state = receiving_dado and done_SI = '1' else -- quando terminarmos de receber�   q   s          n      next_state <= receiving_dado when present_state = initial and serial_in = '0' else -- recebe o start bit�   a   c          Y      type state_type is (initial, receiving_dado, calculando, transmitindo_dado, ended);�   O   Q          4        haso: out bit_vector(255 downto 0); --- dado�   N   P        4        msgi: in bit_vector(511 downto 0);  --- dado5��    N   0                 	                    �    O   0                 ;	                    �    a   -                 2                    �    a   N                 S                    �    q                    �                    �    r   >                 j                    �    s                    �                    �    s   n                                     �    t   !                 Q                    �    u   <                 �                    �    v                    E                    �    {   8                 ,                    �    }   8                 �                    �    �                    �                    �    �   F                 "                    �    Q  A                 0                    �    Q  M                 �0                    �    _  G                 {4                    �    `  C                 �4                    �    b                   J5                    �    d                   �5                    �    e                   6                    5�_�                     �        ����                                                                                                                                                                                                                                                                                                                                                             f)FF    �   �   �          3        contagem_unsigned <= contagem_unsigned + 1;�   �   �          )        --   contagem_unsigned <= "0000";�   �   �          &          contagem_unsigned <= "0000";�   �   �          .        elsif contagem_unsigned=(WIDTH+1) then�   �   �          M          serial_o <= data(to_integer(contagem_unsigned)-1); --saindo datatas�   �   �          L        elsif ((contagem_unsigned > 0) and (contagem_unsigned<WIDTH+1)) then�   �   �          #        if contagem_unsigned=0 then�   �   �          $        contagem_unsigned <= "0000";�   �   �          3    signal contagem_unsigned: unsigned(3 downto 0);�   �   �        ,    signal contagem: bit_vector(3 downto 0);5��    �                    �                    �    �                                        �    �                    �                     �    �                    /!                    �    �                    �!                    �    �   ,                 �!                    �    �   &                 �!                    �    �                    4"                    �    �   
                 �"                    �    �                    v#                    �    �                    �#                    �    �                    �#                    5�_�                    O        ����                                                                                                                                                                                                                                                                                                                                                             f)F     �   N   P        4        msgi: in bit_vector(511 downto 0);  --- data�   O   Q          4        haso: out bit_vector(255 downto 0); --- data�   a   c          Y      type state_type is (initial, receiving_data, calculando, transmitindo_data, ended);�   q   s          n      next_state <= receiving_data when present_state = initial and serial_in = '0' else -- recebe o start bit�   r   t          z                    calculando when present_state = receiving_data and done_SI = '1' else -- quando terminarmos de receber�   s   u          �                    receiving_data when present_state = calculando and serial_in = '0' else -- receiving um data no meio do caculo�   t   v          ~                    transmitindo_data when present_state = calculando and done_MS = '1' else -- quando terminarmos de calcular�   u   w          s                    ended when present_state = transmitindo_data and done_SO = '1' else -- terminamos de trasnmitir�   v   x          Z                    receiving_data when present_state = ended and serial_in = '0'; -- loop�   {   }          A      reset_SO <= '0' when present_state = transmitindo_data else�   }             A      start_SO <= '1' when present_state = transmitindo_data else�   �   �          .    signal data: bit_vector(WIDTH-1 downto 0);�   �   �          K          serial_o <= data(to_integer(contagem_unsigned)-1); --saindo datas�  Q  S          s    signal serial_sig, shift_sig, zero_sig, enable_sig, bit_sig, data_sig, data_sig_stop, clr10_sig, clr4_sig: bit;�  _  a          Z                  waiting_stop_bits when present_state = receiving and data_sig = '1' else�  `  b          [                  ended when present_state = waiting_stop_bits and data_sig_stop = '1' else�  b  d               -- Setting datas de controle�  d  f          q    data_sig <= counter10_out(3) and not(counter10_out(2)) and counter10_out(1) and not(counter10_out(0)); --1010�  e  g          v    data_sig_stop <= counter10_out(3) and counter10_out(2) and not(counter10_out(1)) and not(counter10_out(0)); --11005��    N   0                 	                    �    O   0                 9	                    �    a   -                 .                    �    a   L                 M                    �    q                    �                    �    r   >                 `                    �    s                    �                    �    s   l                 	                    �    t   !                 A                    �    u   <                 �                    �    v                    1                    �    {   8                                     �    }   8                 o                    �    �                    �                    �    �   F                 "                    �    Q  A                 a0                    �    Q  K                 k0                    �    _  G                 Y4                    �    `  C                 �4                    �    b                   $5                    �    d                   p5                    �    e                   �5                    5�_�                    b        ����                                                                                                                                                                                                                                                                                                                                                             f)E�     �   a   c        W      type state_type is (initial, receiving_dado, calculando, transmitindo_dado, end);�   u   w          q                    end when present_state = transmitindo_dado and done_SO = '1' else -- terminamos de trasnmitir�   v   x          X                    receiving_dado when present_state = end and serial_in = '0'; -- loop�  P  R          R    type state_type is (initial, waiting_zero, receiving, waiting_stop_bits, end);�  V  X          k    signal state_initial, state_waiting_zero, state_receiving, state_end, tick: bit; -- sinais para debugar�  a  c          Y                  end when present_state = waiting_stop_bits and dado_sig_stop = '1' else�  b  d          I                  waiting_zero when present_state = end and start = '1'; �  j  l          2    clr10_sig <= '1' when present_state = end else�  u  w          L    parity_bit <= registrador_out((WIDTH + 1) - 1) when present_state = end;�  v  x          2    done <= '1' when present_state = end else '0';�  |  ~          7    state_end <= '1' when present_state = end else '0';5��    a   R                 S                    �    u                    �                    �    v   8                 G                    �    P  M                 �/                    �    V  E                 �1                    �    a                   �4                    �    b  4                 5                    �    j  *                 �7                    �    u  H                 ,;                    �    v  %                 V;                    �    |  
                 �<                    �    |  *                 �<                    5�_�                   {   !    ����                                                                                                                                                                                                                                                                                                                                                             f)Ec     �  z  |        N    estado_esperando_zero <= '1' /hen present_state = esperando_zero else '0';5��    z  !                 I<                    5�_�              
   	  t   /    ����                                                                                                                                                                                                                                                                                                                                                             f)EE     �  s  u        h    CONTADOR10C: counter generic map(WIDTH => 4 port map(bit_sig, clr10_sig, enable_sig, counter10_out);5��    s  /                  �:                     5�_�                   r   N    ����                                                                                                                                                                                                                                                                                                                                                             f)E2     �  q  s        �    REGISTERC: registrador_serial_input generic map(TAMANHO_REG => (WIDTH + 1) port map(shift_sig, serial_data, registrador_out);5��    q  N                  �9                     5�_�                   r   Q    ����                                                                                                                                                                                                                                                                                                                                                             f)E!     �  q  s        �    REGISTRADORC: registrador_serial_input generic map(TAMANHO_REG => (WIDTH + 1) port map(shift_sig, serial_data, registrador_out);5��    q  Q                  �9                     5�_�                             ����                                                                                                                                                                                                                                                                                                                                                             f)D�     �                  entity clock_divider is�   	                 end clock_divider;�                (    architecture arc of clock_divider is�   S   U          $      -- component clock_divider4 is�   Y   [                 component clock_divider is�   �   �          ?      clockTransmissao: clock_divider port map(clock, '0', CT);�   �   �          @      -- clockRecepcao: clock_divider4 port map(clock, '0', CR);5��                        X                     �    	                    �                     �                        	                    �    S                    �	                    �    Y                    .
                    �    �                                        �    �                    N                    5��