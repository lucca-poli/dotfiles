Vim�UnDo� �������0it��F�7��t���S8�	�   �                  	       	   	   	    f=    _�                     �        ����                                                                                                                                                                                                                                                                                                                            �         
          V       f=X     �   �   �       I   entity ch is   
    port (   2        x , y , z : in bit_vector (31 downto 0 ) ;   (        q : out bit_vector (31 downto 0)       ) ;       end ch;          #    architecture ch_arch of ch is             begin   /            q <= (x and y) xor ((not x) and z);       end architecture;              entity sum0 is   
    port (   *        x : in bit_vector (31 downto 0 ) ;   (        q : out bit_vector (31 downto 0)       ) ;       end sum0;          '    architecture sum0_arch of sum0 is             begin   9            q <= (x ror 2) xor (x ror 13) xor (x ror 22);       end architecture;              entity sum1 is   
    port (   *        x : in bit_vector (31 downto 0 ) ;   (        q : out bit_vector (31 downto 0)       ) ;       end sum1;          '    architecture sum1_arch of sum1 is             begin   :            q <=  (x ror 6) xor (x ror 11) xor (x ror 25);       end architecture;              entity maj is   
    port (   2        x , y , z : in bit_vector (31 downto 0 ) ;   (        q : out bit_vector (31 downto 0)       );       end maj ;          %    architecture maj_arch of maj is             begin   7            q <= (x and y) xor (x and z) xor (y and z);       end architecture;              entity sigma0 is   
    port (   *        x : in bit_vector (31 downto 0 ) ;   (        q : out bit_vector (31 downto 0)       ) ;       end sigma0 ;          +    architecture sigma0_arch of sigma0 is             begin   8            q <= (x ror 7) xor (x ror 18) xor (x srl 3);       end architecture;              entity sigma1 is   
    port (   *        x : in bit_vector (31 downto 0 ) ;   (        q : out bit_vector (31 downto 0)       ) ;       end sigma1;          +    architecture sigma1_arch of sigma1 is             begin   :            q <= (x ror 17) xor (x ror 19) xor (x srl 10);       end architecture;           5��    �       I               7      �              5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f=Y    �   �   �           5��    �                      7                     5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �         R          V       f=�     �   �   �       ]   entity stepfun is   port (   M        ai , bi , ci , di , ei , fi , gi , hi : in bit_vector (31 downto 0 );   *        kpw : in bit_vector (31 downto 0);   L        ao , bo , co , do , eo , fo , go , ho : out bit_vector (31 downto 0)       );   end stepfun ;       &architecture stepfunarch of stepfun is       component ch is           port (   1            x, y, z: in bit_vector (31 downto 0);   +            q: out bit_vector (31 downto 0)   
        );       end component;           component maj is            port (   1            x, y, z: in bit_vector (31 downto 0);   +            q: out bit_vector (31 downto 0)   
        );       end component;           component sum0 is            port (   ,            x : in bit_vector (31 downto 0);   ,            q : out bit_vector (31 downto 0)               );       end component;           component sum1 is           port (   +            x: in bit_vector (31 downto 0);   +            q: out bit_vector (31 downto 0)   
        );       end component;           component sigma0 is           port (   +            x: in bit_vector (31 downto 0);   +            q: out bit_vector (31 downto 0)   
        );       end component;           component sigma1 is           port (   +            x: in bit_vector (31 downto 0);   +            q: out bit_vector (31 downto 0)   
        );       end component;           component adder32 is           port (   .            x, y: in  bit_vector(31 downto 0);   +            q: out  bit_vector(31 downto 0)   
        );       end component;          '    signal s1: bit_vector(31 downto 0);   '    signal s2: bit_vector(31 downto 0);   '    signal s3: bit_vector(31 downto 0);   '    signal s4: bit_vector(31 downto 0);   '    signal s5: bit_vector(31 downto 0);   '    signal s6: bit_vector(31 downto 0);       )    signal ch_s: bit_vector(31 downto 0);   *    signal maj_s: bit_vector(31 downto 0);   +    signal sum0_s: bit_vector(31 downto 0);   +    signal sum1_s: bit_vector(31 downto 0);       	    begin   )        sSUM0: sum0 port map(ai, sum0_s);   *        sSUM1: sum1 port map (ei, sum1_s);   ,        sCH: ch port map (ei, fi, gi, ch_s);   .        sMAJ: maj port map(ai, bi, ci, maj_s);              .        PSOMA1: adder32 port map(hi, kpw, s1);   /        PSOMA2: adder32 port map(ch_s, s1, s2);   1        PSOMA3: adder32 port map(sum1_s, s2, s3);   -        PSOMA4: adder32 port map(di, s3, s4);   0        PSOMA5: adder32 port map(maj_s, s3, s5);   1        PSOMA6: adder32 port map(sum0_s, s5, s6);               ao <= s6;           bo <= ai;           co <= bi;           do <= ci;           eo <= s4;           fo <= ei;           go <= fi;           ho <= gi;              end architecture;5��    �       ]               �&      �	              5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f=�    �   �   �           5��    �                      �&                     5�_�      	             �        ����                                                                                                                                                                                                                                                                                                                            �          �           V       f=     �   �   �       4   entity adder32 is   
    port (   *        x, y: in  bit_vector(31 downto 0);   '        q: out  bit_vector(31 downto 0)       );   end entity adder32;       $architecture Archadder of adder32 is       component soma is           port (                a, b, carry: in bit;               sum, cout: out bit   
        );       end component;       (    signal aux: bit_vector(31 downto 0);   begin   9    SOMA0:  soma port map(x(0), y(0), '0', q(0), aux(0));   <    SOMA1:  soma port map(x(1), y(1), aux(0), q(1), aux(1));   <    SOMA2:  soma port map(x(2), y(2), aux(1), q(2), aux(2));   <    SOMA3:  soma port map(x(3), y(3), aux(2), q(3), aux(3));   <    SOMA4:  soma port map(x(4), y(4), aux(3), q(4), aux(4));   <    SOMA5:  soma port map(x(5), y(5), aux(4), q(5), aux(5));   <    SOMA6:  soma port map(x(6), y(6), aux(5), q(6), aux(6));   <    SOMA7:  soma port map(x(7), y(7), aux(6), q(7), aux(7));   <    SOMA8:  soma port map(x(8), y(8), aux(7), q(8), aux(8));   <    SOMA9:  soma port map(x(9), y(9), aux(8), q(9), aux(9));   @    SOMA10: soma port map(x(10), y(10), aux(9), q(10), aux(10));   A    SOMA11: soma port map(x(11), y(11), aux(10), q(11), aux(11));   A    SOMA12: soma port map(x(12), y(12), aux(11), q(12), aux(12));   A    SOMA13: soma port map(x(13), y(13), aux(12), q(13), aux(13));   A    SOMA14: soma port map(x(14), y(14), aux(13), q(14), aux(14));   A    SOMA15: soma port map(x(15), y(15), aux(14), q(15), aux(15));   A    SOMA16: soma port map(x(16), y(16), aux(15), q(16), aux(16));   A    SOMA17: soma port map(x(17), y(17), aux(16), q(17), aux(17));   A    SOMA18: soma port map(x(18), y(18), aux(17), q(18), aux(18));   A    SOMA19: soma port map(x(19), y(19), aux(18), q(19), aux(19));   A    SOMA20: soma port map(x(20), y(20), aux(19), q(20), aux(20));   A    SOMA21: soma port map(x(21), y(21), aux(20), q(21), aux(21));   A    SOMA22: soma port map(x(22), y(22), aux(21), q(22), aux(22));   A    SOMA23: soma port map(x(23), y(23), aux(22), q(23), aux(23));   A    SOMA24: soma port map(x(24), y(24), aux(23), q(24), aux(24));   A    SOMA25: soma port map(x(25), y(25), aux(24), q(25), aux(25));   A    SOMA26: soma port map(x(26), y(26), aux(25), q(26), aux(26));   A    SOMA27: soma port map(x(27), y(27), aux(26), q(27), aux(27));   A    SOMA28: soma port map(x(28), y(28), aux(27), q(28), aux(28));   A    SOMA29: soma port map(x(29), y(29), aux(28), q(29), aux(29));   A    SOMA30: soma port map(x(30), y(30), aux(29), q(30), aux(30));   A    SOMA31: soma port map(x(31), y(31), aux(30), q(31), aux(31));       end architecture Archadder;    5��    �       4               7      �	              5�_�                  	   �        ����                                                                                                                                                                                                                                                                                                                            �          �           V       f=    �   �   �           5��    �                      6                     5�_�                   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        f=�     �      �        5��           u               �      !              5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        f=�     �   ~   �        5��    ~                      �                     5�_�                             ����                                                                                                                                                                                                                                                                                                                                                  V        f=�    �   ~   �        5��    ~                      �                     5��