Vim�UnDo� It}�o�d_�����I�<�����i�57���   @          '         �       �   �   �    fB��    _�                         !    ����                                                                                                                                                                                                                                                                                                                                                             f�    �      !   ?      #	constant test_size: positive := 4;5��       !                                     5�_�                   7   
    ����                                                                                                                                                                                                                                                                                                                            7          7   
       v       f��    �   6   8   ?      			assert check = asserts(i)5��    6   
                 �                    5�_�                   7   
    ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f�_     �   6   8   ?      			assert false5��    6   
                 �                    5�_�      	              7       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f�e     �   6   8   ?      			assert check = asserts5��    6                     �                     5�_�      
           	   7       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f�e     �   6   8   ?      			assert check = asserts()5��    6                     �                     5�_�   	              
   9       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f�y     �   9   ;   ?    �   9   :   ?    5��    9                      q              �       5�_�   
                 :       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f��     �   9   ;   @      �				report "Entrada: " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    9                    }                    �    9                    �                    5�_�                    :       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f��     �   9   ;   @      �				report "haso0 : " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    9                     �                     5�_�                    :   ,    ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f��     �   9   ;   @      �				report "haso0: " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    9   ,                 �                    5�_�                    :   8    ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f��     �   9   ;   @      �				report "haso0: " &  to_hstring(unsigned(check)) & " Esperado: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    9   8                 �                    5�_�                    :   ^    ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f��     �   9   ;   @      �				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    9   ^                 �                    5�_�                    :   h    ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f��     �   9   ;   @      �				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada: " & to_hstring(unsigned(datas(i))) & " Recebido: " & to_hstring(unsigned(check))5��    9   h       .           �      .               5�_�                    :   h    ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f��     �   9   ;   @      h				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada: " & to_hstring(unsigned(datas(i)))5��    9   h                  �                     5�_�                    ;       ����                                                                                                                                                                                                                                                                                                                            :   h       7          V   t    f��    �   ;   @   @    �   ;   <   @    5��    ;                      �              4      5�_�                    ?   D    ����                                                                                                                                                                                                                                                                                                                            :   h       7          V   t    f��    �   >   @   D      i				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada: " & to_hstring(unsigned(datas(i)));5��    >   D                                       5�_�                    4       ����                                                                                                                                                                                                                                                                                                                                                             f
�     �   3   5   D      			wait for 4*half_period;5��    3                    h                    5�_�                    ;       ����                                                                                                                                                                                                                                                                                                                                                             f
�    �   :   <   D      			wait for 4*half_period;5��    :                    �                    5�_�                    !   =    ����                                                                                                                                                                                                                                                                                                                            !   7       !   <       v   ?    fK     �       "   D      L	constant datas: ByteArray(test_size - 1 downto 0) := (x"00", x"01", x"02");5��        =                  Q                     5�_�                    !   =    ����                                                                                                                                                                                                                                                                                                                            !   7       !   <       v   ?    fK     �       "   D      M	constant datas: ByteArray(test_size - 1 downto 0) := (x"00",  x"01", x"02");�   !   "   D    5��        >                  R                     5�_�                   "   F    ����                                                                                                                                                                                                                                                                                                                            "   F       "   :       v   =    fU    �   !   #   D      a	constant asserts: DwordArray(test_size - 1 downto 0) := (x"DA5698BE", x"B8A4E897", x"27D75F9C");�   "   #   D    5��    !   G                  �                     5�_�                        "    ����                                                                                                                                                                                                                                                                                                                            "   F       "   :       v   =    fd    �      !   D      #	constant test_size: positive := 3;5��       !                                     5�_�                   !   >    ����                                                                                                                                                                                                                                                                                                                            !   >       !   D       v   G    fV     �       "   D      S	constant datas: ByteArray(test_size - 1 downto 0) := (x"00", x"00", x"01", x"02");5��        >                  R                     5�_�                   !   D    ����                                                                                                                                                                                                                                                                                                                            !   >       !   D       v   G    fY     �       "   D      L	constant datas: ByteArray(test_size - 1 downto 0) := (x"00", x"01", x"02");�   !   "   D    5��        E                  Y                     5�_�                     "   F    ����                                                                                                                                                                                                                                                                                                                            "   F       "   R       v   U    fj     �   !   #   D      n	constant asserts: DwordArray(test_size - 1 downto 0) := (x"DA5698BE", x"DA5698BE", x"B8A4E897", x"27D75F9C");5��    !   F                  �                     5�_�      H               "   R    ����                                                                                                                                                                                                                                                                                                                                                             fl    �   !   #   D      a	constant asserts: DwordArray(test_size - 1 downto 0) := (x"DA5698BE", x"B8A4E897", x"27D75F9C");�   "   #   D    5��    !   S                  �                     5�_�       I   !       H   #   	    ����                                                                                                                                                                                                                                                                                                                                                             f=     �   #   %   E          �   #   %   D    5��    #                      �                     �    #                                          �    #                                        �    #                                          �    #                                          �    #                                        �    #                                          �    #                                          �    #                 
                
       �    #                                          �    #                                          �    #                                          �    #                                          �    #                                          �    #                                          �    #                                          �    #                                          �    #                                          �    #                 
                
       �    #          
                
              �    #                 
                
       5�_�   H   J           I   $       ����                                                                                                                                                                                                                                                                                                                                                             f=     �   #   %   E          constant exp8: bit_vector5��    #                                          5�_�   I   K           J   $       ����                                                                                                                                                                                                                                                                                                                                                             f=     �   #   %   E          constant exp8: bit_vector()5��    #                                          5�_�   J   O           K   $   +    ����                                                                                                                                                                                                                                                                                                                                                             f=     �   #   %   E      +    constant exp8: bit_vector(511 downto 0)5��    #   +                  (                     �    #   +                 (                    5�_�   K   P   M       O   $   /    ����                                                                                                                                                                                                                                                                                                                                                             f='     �   #   %   E      0    constant exp8: bit_vector(511 downto 0) := ;5��    #   /                  ,                     5�_�   O   Q           P   $   0    ����                                                                                                                                                                                                                                                                                                                                                             f='     �   #   %   E      1    constant exp8: bit_vector(511 downto 0) := x;5��    #   0                  -                     5�_�   P   R           Q   $   1    ����                                                                                                                                                                                                                                                                                                                                                             f=)     �   #   %   E      3    constant exp8: bit_vector(511 downto 0) := x"";�   $   %   E    5��    #   1               @   .              @       5�_�   Q   S           R   $   1    ����                                                                                                                                                                                                                                                                                                                                                             f=I     �   $   %   F      ";�   #   &   E      s    constant exp8: bit_vector(511 downto 0) := x"0f2c074831ecb6102001c11062fd0e5b92b5addd37fa5dca05209e48e21a3845";�   $   %   E    5��    #   1       @           .      @               �    #   1                  .              �       �    #   �                  �                     5�_�   R   T           S   $   �    ����                                                                                                                                                                                                                                                                                                                                                             f=S     �   $   &   E    �   $   %   E    5��    $                      �              �       5�_�   S   U           T   %       ����                                                                                                                                                                                                                                                                                                                                                             f=Z     �   $   &   F      �    constant exp8: bit_vector(511 downto 0) := x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333";5��    $                  	   �              	       5�_�   T   W           U   %   :    ����                                                                                                                                                                                                                                                                                                                                                             f=�     �   $   &   F      �    constant exp8_expected: bit_vector(511 downto 0) := x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333";5��    $   :       �           �      �               5�_�   U   X   V       W   %   :    ����                                                                                                                                                                                                                                                                                                                                                             f=�     �   %   &   G      ";�   $   '   F      <    constant exp8_expected: bit_vector(511 downto 0) := x"";�   %   &   F    5��    $   :                  �              A       �    $   z                  +                     5�_�   W   \           X   *   1    ����                                                                                                                                                                                                                                                                                                                            +   8       *   2       V   y    f=�     �   )   ,   F      2	Qword <= data&data&data&data&data&data&data&data;   9	msgi <= Qword&Qword&Qword&Qword&Qword&Qword&Qword&Qword;5��    )                     x      m       s       5�_�   X   ]   Y       \   3   %    ����                                                                                                                                                                                                                                                                                                                            +   8       *   2       V   y    f=�     �   2   4   F      &		for i in test_size - 1 downto 0 loop5��    2                     \      '       *       5�_�   \   ^           ]   5       ����                                                                                                                                                                                                                                                                                                                            +   8       *   2       V   y    f=�     �   4   6   F      			data <= datas(i);5��    4                     �                    5�_�   ]   _           ^   B   
    ����                                                                                                                                                                                                                                                                                                                            +   8       *   2       V   y    f=�     �   A   C   F      		end loop;5��    A                     |	                    5�_�   ^   `           _   ,       ����                                                                                                                                                                                                                                                                                                                            +   8       *   2       V   y    f=�     �   +   -   F      	check <= haso(31 downto 0);5��    +                     �                     5�_�   _   a           `   9       ����                                                                                                                                                                                                                                                                                                                            9          9          v   $    f=	     �   8   :   F      			assert check = asserts(i)5��    8          
          �      
              �    8                                           �    8                     �                     �    8                    �                    �    8                    �                    �    8                    �                    �    8                    �                    5�_�   `   b           a   >       ����                                                                                                                                                                                                                                                                                                                            9          9          v   $    f=     �   =   ?   F      			assert check = asserts(i)5��    =          
          Q      
              �    =                     S                     �    =                     R                     �    =                    Q                    �    =                    Q                    �    =                    Q                    5�_�   a   c           b   :   .    ����                                                                                                                                                                                                                                                                                                                            :   .       :   5       v   A    f=;     �   9   ;   F      �				report "Entrada: " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    9   .                 :                    �    9   .                 :                    �    9   .                 :                    �    9   .                 :                    �    9   .                 :                    �    9   .                 :                    5�_�   b   d           c   ?   .    ����                                                                                                                                                                                                                                                                                                                            :   .       :   5       v   A    f=K     �   >   @   F      �				report "Entrada: " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    >   .                 �                    �    >   .                 �                    �    >   .                 �                    �    >   .                 �                    5�_�   c   e           d   :   [    ����                                                                                                                                                                                                                                                                                                                            :   .       :   5       v   A    f=T     �   9   ;   F      �				report "Entrada: " &  to_hstring(unsigned(exp8)) & " Esperado: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    9   [       
          g      
              �    9   [                 g                    �    9   [                 g                    �    9   [                 g                    �    9   [                 g                    �    9   [                 g                    5�_�   d   f           e   ?   [    ����                                                                                                                                                                                                                                                                                                                            :   .       :   5       v   A    f=h     �   >   @   F      �				report "Entrada: " &  to_hstring(unsigned(exp8)) & " Esperado: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    >   [       
          �      
              �    >   [                 �                    �    >   [                 �                    �    >   [                 �                    �    >   [                 �                    5�_�   e   g           f   <   ^    ����                                                                                                                                                                                                                                                                                                                            :   .       :   5       v   A    f=r     �   ;   =   F      i				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada: " & to_hstring(unsigned(datas(i)));5��    ;   ^                                     �    ;   ^                                     �    ;   ^                                     �    ;   ^                                     �    ;   ^                                     �    ;   ^                                     5�_�   f   h           g   A   ]    ����                                                                                                                                                                                                                                                                                                                            :   .       :   5       v   A    f={    �   @   B   F      h				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada " & to_hstring(unsigned(datas(i)));5��    @   ]                 c	                    �    @   ]                 c	                    �    @   ]                 c	                    �    @   ]                 c	                    5�_�   g   i           h          ����                                                                                                                                                                                                                                                                                                                            :   .       :   5       v   A    f=�    �         F      '	signal check: bit_vector(31 downto 0);5��                        '                    5�_�   h   j           i   %   '    ����                                                                                                                                                                                                                                                                                                                            :   .       :   5       v   A    f=�    �   $   &   F      |    constant exp8_expected: bit_vector(511 downto 0) := x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd";5��    $   '                 �                    5�_�   i   k           j   *        ����                                                                                                                                                                                                                                                                                                                                                             fBw�     �               F   library ieee;   use ieee.numeric_bit.all;   use std.textio.all;       entity dut is end;       architecture dut_arch of dut is       	component multisteps is   		port (clk, rst : in  bit;   ,				msgi     : in  bit_vector(511 downto 0);   )				haso		: out bit_vector(255 downto 0);   				done		: out bit   		);   	end component multisteps;           	signal clk: bit := '0';   	signal rst: bit := '0';   	signal done: bit;   	signal finished: bit := '0';   %	signal data: bit_vector(7 downto 0);   '	signal Qword: bit_vector(63 downto 0);   '	signal msgi: bit_vector(511 downto 0);   (	signal check: bit_vector(255 downto 0);   '	signal haso: bit_vector(255 downto 0);       F	type ByteArray is array (natural range <>) of bit_vector(7 downto 0);   H	type DwordArray is array (natural range <>) of bit_vector(31 downto 0);           #	constant test_size: positive := 4;   S	constant datas: ByteArray(test_size - 1 downto 0) := (x"00", x"01", x"00", x"02");   n	constant asserts: DwordArray(test_size - 1 downto 0) := (x"DA5698BE", x"B8A4E897", x"DA5698BE", x"27D75F9C");   %	constant half_period : time := 1 ns;   �    constant exp8: bit_vector(511 downto 0) := x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333";   |    constant exp8_expected: bit_vector(255 downto 0) := x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd";   	   begin       @	clk <= not clk after half_period when finished /= '1' else '0';   5	-- Qword <= data&data&data&data&data&data&data&data;   <	-- msgi <= Qword&Qword&Qword&Qword&Qword&Qword&Qword&Qword;   	check <= haso;       	exp4dut: multisteps   '	port map(clk, rst, msgi, haso,  done);   	   	st: process   	begin   )		-- for i in test_size - 1 downto 0 loop   			rst <= '1';   			-- data <= datas(i);   			wait for 16*half_period;   			rst <= '0';    			wait until rising_edge(done);   			assert check = exp8_expected   �				report "Entrada: " &  to_hstring(unsigned(exp8)) & " Esperado: " & to_hstring(unsigned(exp8_expected)) & " Recebido: " & to_hstring(unsigned(check))   				severity note;   e				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada: " & to_hstring(unsigned(exp8));   			wait for 31*half_period;   			assert check = exp8_expected   �				report "Entrada: " &  to_hstring(unsigned(exp8)) & " Esperado: " & to_hstring(unsigned(exp8_expected)) & " Recebido: " & to_hstring(unsigned(check))   				severity note;   d				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada " & to_hstring(unsigned(exp8));   		-- end loop;   		finished <= '1';   		wait;   	end process;   end;5�5�_�   j   l           k   $       ����                                                                                                                                                                                                                                                                                                                                                             fBw�     �   $   &   F    �   $   %   F    5��    $                      �              �       5�_�   k   m           l   $       ����                                                                                                                                                                                                                                                                                                                                                             fBw�     �   #   %   G      �    constant exp8: bit_vector(511 downto 0) := x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333";5��    #                                        5�_�   l   n           m       !    ����                                                                                                                                                                                                                                                                                                                                                             fBx     �      !   G      #	constant test_size: positive := 4;5��       !                                     5�_�   m   o           n   $       ����                                                                                                                                                                                                                                                                                                                            $          $   +       v   +    fBx     �   #   %   G      �    constant datas: bit_vector(511 downto 0) := x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333";5��    #                                        �    #                                        �    #                                          �    #                                        5�_�   n   p           o   $       ����                                                                                                                                                                                                                                                                                                                            $          $   +       v   +    fBxM     �   #   %   G      �    constant datas: InArray := x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333";5��    #                                          5�_�   o   q           p   $       ����                                                                                                                                                                                                                                                                                                                            $          $   +       v   +    fBxN     �   #   %   G      �    constant datas: InArray() := x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333";5��    #                                          �    #                 	                	       �    #          	                	              �    #                                        �    #   (                  (                     �    #   '                 '                    �    #   *                 *                    �    #   *                 *                    �    #   *                 *                    5�_�   p   r           q          ����                                                                                                                                                                                                                                                                                                                            $          $   +       v   +    fBxX     �         G      F	type ByteArray is array (natural range <>) of bit_vector(7 downto 0);5��              	          e      	              �                        e                    �                        e                    �                        e                    5�_�   q   s           r      9    ����                                                                                                                                                                                                                                                                                                                            $          $   +       v   +    fBx^     �         G      D	type InArray is array (natural range <>) of bit_vector(7 downto 0);5��       8                 �                    �       8                 �                    5�_�   r   t           s      ;    ����                                                                                                                                                                                                                                                                                                                            $          $   +       v   +    fBxc     �         G      H	type DwordArray is array (natural range <>) of bit_vector(31 downto 0);5��       ;                 �                    5�_�   s   u           t          ����                                                                                                                                                                                                                                                                                                                            $          $   +       v   +    fBxh     �         G      I	type DwordArray is array (natural range <>) of bit_vector(255 downto 0);5��              
          �      
              �                         �                     �                         �                     �                        �                    �                         �                     �                         �                     �       
                  �                     �       	                  �                     �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    5�_�   t   v           u          ����                                                                                                                                                                                                                                                                                                                            $          $   +       v   +    fBxn     �         G      F	type InArray is array (natural range <>) of bit_vector(255 downto 0);5��                        �                    5�_�   u   w           v       !    ����                                                                                                                                                                                                                                                                                                                            $          $   +       v   +    fBxt     �      !   G      %	constant test_size: positive := 512;5��       !                                     5�_�   v   x           w   &       ����                                                                                                                                                                                                                                                                                                                            $          $   +       v   +    fBx�     �   %   '   G      |    constant exp8_expected: bit_vector(255 downto 0) := x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd";5��    %                    z                    �    %                    z                    �    %                                          �    %                     ~                     �    %                     }                     �    %                     |                     �    %                     {                     �    %                    z                    �    %                    z                    �    %                    z                    �    %                    z                    5�_�   w   y           x   &       ����                                                                                                                                                                                                                                                                                                                            &          &          v       fBx�     �   %   '   G      v    constant asserts: bit_vector(255 downto 0) := x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd";5��    %          
           �      
               5�_�   x   z           y   &       ����                                                                                                                                                                                                                                                                                                                            &          &          v       fBx�     �   %   '   G      l    constant asserts: (255 downto 0) := x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd";5��    %                     �                     5�_�   y   {           z   &       ����                                                                                                                                                                                                                                                                                                                            &          &          v       fBx�     �   %   '   G      ^    constant asserts:  := x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd";5��    %                     �                     �    %                     �                     �    %                     �                     �    %                    �                    �    %                    �                    �    %                    �                    5�_�   z   |           {   &       ����                                                                                                                                                                                                                                                                                                                            &          &          v       fBx�     �   %   '   G      f    constant asserts: OutArray := x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd";5��    %                     �                     5�_�   {   }           |   &       ����                                                                                                                                                                                                                                                                                                                            &          &          v       fBx�     �   %   '   G      h    constant asserts: OutArray() := x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd";5��    %                     �                     �    %   !                  �                     �    %                      �                     �    %                 	   �             	       �    %          	          �      	              �    %                    �                    �    %   -                 �                    �    %   -                 �                    �    %   -                 �                    5�_�   |   ~           }   &   :    ����                                                                                                                                                                                                                                                                                                                            &          &          v       fBx�     �   %   '   G      ~    constant asserts: OutArray(test_size - 1 downto 0) := x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd";5��    %   :                  �                     5�_�   }              ~   &   ;    ����                                                                                                                                                                                                                                                                                                                            &          &          v       fBx�     �   %   '   G          constant asserts: OutArray(test_size - 1 downto 0) := (x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd";5��    %                     m      �       �       5�_�   ~   �              %   }    ����                                                                                                                                                                                                                                                                                                                            &          &          v       fBx�     �   $   %          �    constant exp8: bit_vector(511 downto 0) := x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333";5��    $                      �      �               5�_�      �           �   $   7    ����                                                                                                                                                                                                                                                                                                                            %          %          v       fBx�     �   #   %   F      �    constant datas: InArray(test_size - 1 downto 0) := x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333";5��    #   7                  4                     5�_�   �   �           �   $   8    ����                                                                                                                                                                                                                                                                                                                            %          %          v       fBx�     �   #   %   F      �    constant datas: InArray(test_size - 1 downto 0) := (x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333";5��    #                     �      �       �       5�_�   �   �           �   $   �    ����                                                                                                                                                                                                                                                                                                                            %          %          v       fBx�     �   #   %   F      �    constant datas: InArray(test_size - 1 downto 0) := (x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333");5��    #   �                  �                     �    #   �                 �                    5�_�   �   �           �   $   �    ����                                                                                                                                                                                                                                                                                                                            %          %          v       fBx�     �   #   %   F      �    constant datas: InArray(test_size - 1 downto 0) := (x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333", x);5��    #   �                  �                     5�_�   �   �           �   $   �    ����                                                                                                                                                                                                                                                                                                                            %          %          v       fBx�     �   #   %   F      �    constant datas: InArray(test_size - 1 downto 0) := (x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333", x"");�   $   %   F    5��    #   �                  �                     �    #   �              �   �             �       5�_�   �   �           �   $        ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fBy      �   #   %   F     �    constant datas: InArray(test_size - 1 downto 0) := (x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333", x"4c 61 62 6f 72 61 74 6f 72 69 6f 20 44 69 67 69 74 61 6c 20 65 68 20 6d 75 69 74 6f 20 66 61 63 69 6c 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f 5f");5��    #                      �                     �    #                                          �    #                                          �    #                                          �    #                                           �    #   !                                       �    #   '                  $                     �    #   )                  &                     �    #   +                  (                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #   �                  �                     �    #                     �                     �    #                    �                     �    #                                         �    #                                         �    #                                         �    #   
                                      �    #                    	                     �    #                                         �    #                                         �    #                                         �    #                                         �    #                                         �    #                                         �    #                                         �    #                                         �    #                                         �    #                                          �    #   "                                      �    #   $                 !                     �    #   &                 #                     �    #   (                 %                     �    #   *                 '                     �    #   ,                 )                     �    #   .                 +                     �    #   0                 -                     5�_�   �   �           �   $        ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fBy!     �   #   %   F     5constantdatas:InArray(test_size-1downto0):=(x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333",x"4c61626f7261746f72696f204469676974616c206568206d7569746f20666163696c5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f");5��    #                      �                     5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fBy$     �   #   %   F     9    constantdatas:InArray(test_size-1downto0):=(x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333",x"4c61626f7261746f72696f204469676974616c206568206d7569746f20666163696c5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f");5��    #                     	                     5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fBy&     �   #   %   F     :    constant datas:InArray(test_size-1downto0):=(x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333",x"4c61626f7261746f72696f204469676974616c206568206d7569746f20666163696c5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f");5��    #                                          5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fBy(     �   #   %   F     ;    constant datas :InArray(test_size-1downto0):=(x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333",x"4c61626f7261746f72696f204469676974616c206568206d7569746f20666163696c5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f");5��    #                                          5�_�   �   �           �   $   &    ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fBy,     �   #   %   F     <    constant datas : InArray(test_size-1downto0):=(x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333",x"4c61626f7261746f72696f204469676974616c206568206d7569746f20666163696c5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f");5��    #   &                  #                     5�_�   �   �           �   $   )    ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fBy-     �   #   %   F     =    constant datas : InArray(test_size -1downto0):=(x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333",x"4c61626f7261746f72696f204469676974616c206568206d7569746f20666163696c5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f");5��    #   )                  &                     5�_�   �   �           �   $   (    ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fBy/     �   #   %   F     >    constant datas : InArray(test_size -1 downto0):=(x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333",x"4c61626f7261746f72696f204469676974616c206568206d7569746f20666163696c5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f");5��    #   (                  %                     5�_�   �   �           �   $   1    ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fBy1     �   #   %   F     ?    constant datas : InArray(test_size - 1 downto0):=(x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333",x"4c61626f7261746f72696f204469676974616c206568206d7569746f20666163696c5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f");5��    #   1                  .                     5�_�   �   �           �   $   4    ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fBy3     �   #   %   F     @    constant datas : InArray(test_size - 1 downto 0):=(x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333",x"4c61626f7261746f72696f204469676974616c206568206d7569746f20666163696c5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f");5��    #   4                  1                     5�_�   �   �           �   $   7    ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fBy5     �   #   %   F     A    constant datas : InArray(test_size - 1 downto 0) :=(x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333",x"4c61626f7261746f72696f204469676974616c206568206d7569746f20666163696c5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f");5��    #   7                  4                     5�_�   �   �           �   $   �    ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fBy9     �   #   %   F     B    constant datas : InArray(test_size - 1 downto 0) := (x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333",x"4c61626f7261746f72696f204469676974616c206568206d7569746f20666163696c5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f");5��    #   �                  �                     5�_�   �   �           �   %   ~    ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fByR     �   $   &   F      �    constant asserts: OutArray(test_size - 1 downto 0) := (x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd");5��    $   ~                  �                     5�_�   �   �           �   %   �    ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fByT     �   $   &   F      �    constant asserts: OutArray(test_size - 1 downto 0) := (x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd", x);5��    $   �                  �                     5�_�   �   �           �   %   �    ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fByU     �   $   &   F      �    constant asserts: OutArray(test_size - 1 downto 0) := (x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd", x"");�   %   &   F    5��    $   �               d   �              d       5�_�   �   �           �   %   �    ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fByf     �   $   &   F      �    constant asserts: OutArray(test_size - 1 downto 0) := (x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd", x"29 C1 D0 78 62 F1 52 35 D2 4F F1 2F CD A3 87 EF 49 FF 59 91 B8 57 38 D4 C0 77 22 24 97 65 B8 62");5��    $   �                  �                     5�_�   �   �           �   %   �    ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fByl     �   $   &   F      �    constant asserts: OutArray(test_size - 1 downto 0) := (x"bd02d673ff4e4868c1f015c8ffeb420330b75ee36dbc77d05c6e9b20de7168fd", x"29C1 D0 78 62 F1 52 35 D2 4F F1 2F CD A3 87 EF 49 FF 59 91 B8 57 38 D4 C0 77 22 24 97 65 B8 62");5��    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                  �                     �    $   �                                       5�_�   �   �           �   !   R    ����                                                                                                                                                                                                                                                                                                                            $   �       $  }       v  }    fByt     �       !          S	constant datas: ByteArray(test_size - 1 downto 0) := (x"00", x"01", x"00", x"02");   n	constant asserts: DwordArray(test_size - 1 downto 0) := (x"DA5698BE", x"B8A4E897", x"DA5698BE", x"27D75F9C");5��                                 �               5�_�   �   �           �   7       ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBy|     �   6   8   D      			assert check = exp8_expected5��    6                                          5�_�   �   �           �   3       ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz     �   2   4   D      			-- data <= datas(i);5��    2                     �                    5�_�   �   �           �   1       ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz     �   0   2   D      )		-- for i in test_size - 1 downto 0 loop5��    0                     e      *       '       5�_�   �   �           �   @       ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz     �   ?   A   D      		-- end loop;5��    ?                     n	                    5�_�   �   �           �   7       ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz"     �   6   8   D      			assert check = 5��    6                                          �    6                                        �    6                                        �    6                                        �    6                                        5�_�   �   �           �   7       ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz$     �   6   8   D      			assert check = asserts5��    6                                          5�_�   �   �           �   7       ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz&     �   6   8   D      			assert check = asserts()5��    6                                          5�_�   �   �           �   8   .    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz1     �   7   9   D      �				report "Entrada: " &  to_hstring(unsigned(exp8)) & " Esperado: " & to_hstring(unsigned(exp8_expected)) & " Recebido: " & to_hstring(unsigned(check))5��    7   .                 G                    5�_�   �   �           �   8   3    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz4     �   7   9   D      �				report "Entrada: " &  to_hstring(unsigned(datas)) & " Esperado: " & to_hstring(unsigned(exp8_expected)) & " Recebido: " & to_hstring(unsigned(check))5��    7   3                  L                     5�_�   �   �           �   8   4    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz4     �   7   9   D      �				report "Entrada: " &  to_hstring(unsigned(datas())) & " Esperado: " & to_hstring(unsigned(exp8_expected)) & " Recebido: " & to_hstring(unsigned(check))5��    7   4                  M                     5�_�   �   �           �   8   _    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz8     �   7   9   D      �				report "Entrada: " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(exp8_expected)) & " Recebido: " & to_hstring(unsigned(check))5��    7   _                 x                    �    7   _                 x                    �    7   _                 x                    5�_�   �   �           �   8   f    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz<     �   7   9   D      �				report "Entrada: " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(asserts)) & " Recebido: " & to_hstring(unsigned(check))5��    7   f                                       5�_�   �   �           �   8   g    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz=     �   7   9   D      �				report "Entrada: " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(asserts())) & " Recebido: " & to_hstring(unsigned(check))5��    7   g                  �                     5�_�   �   �           �   :   ^    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBzJ     �   9   ;   D      e				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada: " & to_hstring(unsigned(exp8));5��    9   ^                  $                     5�_�   �   �           �   :   ]    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBzP     �   9   :          a				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada: " & to_hstring(unsigned());5��    9                      �      b               5�_�   �   �           �   <   .    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBzU     �   ;   =   C      �				report "Entrada: " &  to_hstring(unsigned(exp8)) & " Esperado: " & to_hstring(unsigned(exp8_expected)) & " Recebido: " & to_hstring(unsigned(check))5��    ;   .                 0                    �    ;   .                 0                    �    ;   .                 0                    �    ;   .                 0                    �    ;   .                 0                    5�_�   �   �           �   <   3    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBzY     �   ;   =   C      �				report "Entrada: " &  to_hstring(unsigned(datas)) & " Esperado: " & to_hstring(unsigned(exp8_expected)) & " Recebido: " & to_hstring(unsigned(check))5��    ;   3                  5                     5�_�   �   �           �   <   4    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBzZ     �   ;   =   C      �				report "Entrada: " &  to_hstring(unsigned(datas())) & " Esperado: " & to_hstring(unsigned(exp8_expected)) & " Recebido: " & to_hstring(unsigned(check))5��    ;   4                  6                     5�_�   �   �           �   <   _    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz]     �   ;   =   C      �				report "Entrada: " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(exp8_expected)) & " Recebido: " & to_hstring(unsigned(check))5��    ;   _                 a                    �    ;   _                 a                    �    ;   _                 a                    �    ;   _                 a                    �    ;   _                 a                    �    ;   _                 a                    5�_�   �   �           �   <   f    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBzb     �   ;   =   C      �				report "Entrada: " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(asserts)) & " Recebido: " & to_hstring(unsigned(check))5��    ;   f                  h                     5�_�   �   �           �   <   g    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBzb     �   ;   =   C      �				report "Entrada: " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(asserts())) & " Recebido: " & to_hstring(unsigned(check))5��    ;   g                  i                     5�_�   �   �           �   <   �    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBzf     �   ;   =   C      �				report "Entrada: " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    ;   �                 �                    �    ;   �                 �                    �    ;   �                 �                    �    ;   �                 �                    5�_�   �   �           �   >   c    ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBzj    �   =   >          d				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada " & to_hstring(unsigned(exp8));5��    =                      �      e               5�_�   �   �           �   ;       ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz�     �   :   <   B      			assert check = exp8_expected5��    :                    �                    �    :                    �                    �    :                     �                     �    :                     �                     �    :                     �                     �    :                     �                     �    :                     �                     �    :                    �                    �    :                    �                    �    :                    �                    �    :                    �                    5�_�   �   �           �   ;       ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz�     �   :   <   B      			assert check = asserts5��    :                     �                     5�_�   �   �           �   ;       ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fBz�    �   :   <   B      			assert check = asserts()5��    :                     �                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fB{     �         B      %	signal data: bit_vector(7 downto 0);5��                        �                    5�_�   �   �   �       �          ����                                                                                                                                                                                                                                                                                                                            "   �       "  }       v  }    fB{5    �                '	signal Qword: bit_vector(63 downto 0);5��                          �      (               5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            !   �       !  }       v  }    fB{K    �         A      '	signal data: bit_vector(512 downto 0);5��                        �                    5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            !   �       !  }       v  }    fB�    �   &   '          5	-- Qword <= data&data&data&data&data&data&data&data;   <	-- msgi <= Qword&Qword&Qword&Qword&Qword&Qword&Qword&Qword;5��    &                      h      s               5�_�   �               �   '       ����                                                                                                                                                                                                                                                                                                                                                             fB��    �   &   (   @          �   &   (   ?    5��    &                      h                     �    &                     l                     �    &                     m                     �    &                    l                    �    &                    l                    �    &                    l                    5�_�   �       �   �   �          ����                                                                                                                                                                                                                                                                                                                            !   �       !  }       v  }    fB{-     �              5��                          �      (               5�_�   �           �   �          ����                                                                                                                                                                                                                                                                                                                                �          }       v  }    fB{*     �              5��                          �      P               5�_�   X   Z       \   Y   3   %    ����                                                                                                                                                                                                                                                                                                                            +   8       *   2       V   y    f=�     �   2   4        5��    2                      \      '               5�_�   Y   [           Z   A   
    ����                                                                                                                                                                                                                                                                                                                            +   8       *   2       V   y    f=�     �   @   B        5��    @                      O	                     5�_�   Z               [   4       ����                                                                                                                                                                                                                                                                                                                            +   8       *   2       V   y    f=�     �   3   5   D      			-- data <= datas(i);5��    3                     k                    5�_�   U           W   V   %   9    ����                                                                                                                                                                                                                                                                                                                                                             f=�     �   %   &   F    �   $   &   F      �    constant exp8_expected: bit_vector(511 downto 0) := x"000000f8000000000000000000000000000000000000000000000000000000006c204180676974616f204469746f7269626f72612d204c613333352050435333";5��    $   :               �   �              �       5�_�   K   N   L   O   M   $   /    ����                                                                                                                                                                                                                                                                                                                                                             f="     �   $   %   E    �   #   %   E      p    constant exp8: bit_vector(511 downto 0) := 0f2c074831ecb6102001c11062fd0e5b92b5addd37fa5dca05209e48e21a3845;5��    #   /               @   ,              @       5�_�   M               N   $   o    ����                                                                                                                                                                                                                                                                                                                                                             f=$     �   #   %   E      r    constant exp8: bit_vector(511 downto 0) := 0f2c074831ecb6102001c11062fd0e5b92b5addd37fa5dca05209e48e21a3845"";5��    #   o                  l                     5�_�   K           M   L   $   .    ����                                                                                                                                                                                                                                                                                                                                                             f=     �   $   %   E    �   $   %   E  k   library IEEE;   use IEEE.NUMERIC_BIT.all;       entity reg32 is   
    port (   !        rst, clk, enable: in bit;   )        init: in bit_vector(31 downto 0);   &        d: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)       );   end entity reg32;       !architecture Behavior of reg32 is   *    signal value: bit_vector(31 downto 0);   begin              process(rst, clk)   	    begin           if rst = '1' then               value <= init;   4        elsif rising_edge(clk) and enable = '1' then               value <= D;           end if;       end process;           q <= value;          end architecture Behavior;       library IEEE;   use IEEE.NUMERIC_BIT.all;       entity shift_reg512 is   
    port (   !        rst, clk, enable: in bit;   )        data: in bit_vector(31 downto 0);   '        d: in bit_vector(511 downto 0);   '        q: out bit_vector(511 downto 0)       );   end entity shift_reg512;       (architecture Behavior of shift_reg512 is   ,   signal vector: bit_vector(511 downto 0);        begin              process(rst, clk)   	    begin           if rst = '1' then               vector <= d;   4        elsif rising_edge(clk) and enable = '1' then   2            vector <= vector(479 downto 0) & data;           end if;       end process;           q <= vector;          end architecture Behavior;       library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity counter_6bit is   
    port (   C        clk, rst: in bit;                            -- Clock input           done: out bit;   O        count : out unsigned(5 downto 0)       -- 6-bit count output (64 steps)       );   end counter_6bit;       #architecture rtl of counter_6bit is   )    signal counter: unsigned(5 downto 0);       begin              counting: process(clk, rst)   	    begin           if rst = '1' then   '            counter <= (others => '0');               done <= '0';   +        elsif to_integer(counter) = 63 then               done <= '1';   #        elsif rising_edge(clk) then   #            counter <= counter + 1;           end if;       end process counting;           count <= counter;          end architecture rtl;       library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity multisteps is   
    port (           clk, rst : in bit;   +        msgi : in bit_vector(511 downto 0);   ,        haso : out bit_vector(255 downto 0);           done : out bit       );   end multisteps;       !architecture rtl of multisteps is           component stepfun  is           port (   D        	ai, bi, ci, di, ei, fi, gi, hi: in bit_vector(31 downto 0);   ,            kpw: in bit_vector(31 downto 0);   G            ao, bo, co, do, eo, fo, go, ho: out bit_vector(31 downto 0)   
        );       end component;           component reg32 is           port (   %            rst, clk, enable: in bit;   -            init: in bit_vector(31 downto 0);   *            d: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component shift_reg512 is           port (   %            rst, clk, enable: in bit;   -            data: in bit_vector(31 downto 0);   +            d: in bit_vector(511 downto 0);   +            q: out bit_vector(511 downto 0)   
        );       end component;           component counter_6bit  is           port (   G            clk, rst: in bit;                            -- Clock input               done: out bit;   S            count : out unsigned(5 downto 0)       -- 6-bit count output (64 steps)   
        );       end component;           component adder32  is           port (   +            a : in bit_vector(31 downto 0);   +            b : in bit_vector(31 downto 0);   +            s : out bit_vector(31 downto 0)   
        );       end component;           component sigma0 is            port(   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;              component sigma1 is           port(   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           -- Constants   9    constant h0 : bit_vector(31 downto 0) := x"6a09e667";   9    constant h1 : bit_vector(31 downto 0) := x"bb67ae85";   9    constant h2 : bit_vector(31 downto 0) := x"3c6ef372";   9    constant h3 : bit_vector(31 downto 0) := x"a54ff53a";   9    constant h4 : bit_vector(31 downto 0) := x"510e527f";   9    constant h5 : bit_vector(31 downto 0) := x"9b05688c";   9    constant h6 : bit_vector(31 downto 0) := x"1f83d9ab";   9    constant h7 : bit_vector(31 downto 0) := x"5be0cd19";           -- Signals   C    type aux_signals is array (0 to 63) of bit_vector(31 downto 0);        signal k_const: aux_signals;       +    signal iteration: unsigned(5 downto 0);       signal ended: bit;   +    signal w_vec: bit_vector(511 downto 0);   +    signal next_w: bit_vector(31 downto 0);   .    signal current_w: bit_vector(31 downto 0);   .    signal current_k: bit_vector(31 downto 0);   0    signal current_kpw: bit_vector(31 downto 0);       *    signal haso0: bit_vector(31 downto 0);   *    signal haso1: bit_vector(31 downto 0);   *    signal haso2: bit_vector(31 downto 0);   *    signal haso3: bit_vector(31 downto 0);   *    signal haso4: bit_vector(31 downto 0);   *    signal haso5: bit_vector(31 downto 0);   *    signal haso6: bit_vector(31 downto 0);   *    signal haso7: bit_vector(31 downto 0);       7    signal op1, op2, op3, op4: bit_vector(31 downto 0);   '    signal av: bit_vector(31 downto 0);   '    signal bv: bit_vector(31 downto 0);   '    signal cv: bit_vector(31 downto 0);   '    signal dv: bit_vector(31 downto 0);   '    signal ev: bit_vector(31 downto 0);   '    signal fv: bit_vector(31 downto 0);   '    signal gv: bit_vector(31 downto 0);   '    signal hv: bit_vector(31 downto 0);   *    signal a_reg: bit_vector(31 downto 0);   *    signal b_reg: bit_vector(31 downto 0);   *    signal c_reg: bit_vector(31 downto 0);   *    signal d_reg: bit_vector(31 downto 0);   *    signal e_reg: bit_vector(31 downto 0);   *    signal f_reg: bit_vector(31 downto 0);   *    signal g_reg: bit_vector(31 downto 0);   *    signal h_reg: bit_vector(31 downto 0);       begin              -- Assynchronous operations       k_const(0) <= x"428a2f98";       k_const(1) <= x"71374491";       k_const(2) <= x"b5c0fbcf";       k_const(3) <= x"e9b5dba5";       k_const(4) <= x"3956c25b";       k_const(5) <= x"59f111f1";       k_const(6) <= x"923f82a4";       k_const(7) <= x"ab1c5ed5";       k_const(8) <= x"d807aa98";       k_const(9) <= x"12835b01";       k_const(10) <= x"243185be";       k_const(11) <= x"550c7dc3";       k_const(12) <= x"72be5d74";       k_const(13) <= x"80deb1fe";       k_const(14) <= x"9bdc06a7";       k_const(15) <= x"c19bf174";       k_const(16) <= x"e49b69c1";       k_const(17) <= x"efbe4786";       k_const(18) <= x"0fc19dc6";       k_const(19) <= x"240ca1cc";       k_const(20) <= x"2de92c6f";       k_const(21) <= x"4a7484aa";       k_const(22) <= x"5cb0a9dc";       k_const(23) <= x"76f988da";       k_const(24) <= x"983e5152";       k_const(25) <= x"a831c66d";       k_const(26) <= x"b00327c8";       k_const(27) <= x"bf597fc7";       k_const(28) <= x"c6e00bf3";       k_const(29) <= x"d5a79147";       k_const(30) <= x"06ca6351";       k_const(31) <= x"14292967";       k_const(32) <= x"27b70a85";       k_const(33) <= x"2e1b2138";       k_const(34) <= x"4d2c6dfc";       k_const(35) <= x"53380d13";       k_const(36) <= x"650a7354";       k_const(37) <= x"766a0abb";       k_const(38) <= x"81c2c92e";       k_const(39) <= x"92722c85";       k_const(40) <= x"a2bfe8a1";       k_const(41) <= x"a81a664b";       k_const(42) <= x"c24b8b70";       k_const(43) <= x"c76c51a3";       k_const(44) <= x"d192e819";       k_const(45) <= x"d6990624";       k_const(46) <= x"f40e3585";       k_const(47) <= x"106aa070";       k_const(48) <= x"19a4c116";       k_const(49) <= x"1e376c08";       k_const(50) <= x"2748774c";       k_const(51) <= x"34b0bcb5";       k_const(52) <= x"391c0cb3";       k_const(53) <= x"4ed8aa4a";       k_const(54) <= x"5b9cca4f";       k_const(55) <= x"682e6ff3";       k_const(56) <= x"748f82ee";       k_const(57) <= x"78a5636f";       k_const(58) <= x"84c87814";       k_const(59) <= x"8cc70208";       k_const(60) <= x"90befffa";       k_const(61) <= x"a4506ceb";       k_const(62) <= x"bef9a3f7";       k_const(63) <= x"c67178f2";           -- W combinational   <    int1: sigma1 port map(w_vec(63 downto 32), op1); -- t-14   =    int2: sigma0 port map(w_vec(479 downto 448), op2); -- t-1   *    int4: adder32 port map(op1, op2, op3);   [    int3: adder32 port map(w_vec(223 downto 192), w_vec(511 downto 480), op4); -- t-9 and t   -    int5: adder32 port map(op3, op4, next_w);           -- W sequential   L    shf_w: shift_reg512 port map (rst, clk, not ended, next_w, msgi, w_vec);       B    get_kpw: adder32 port map (current_w, current_k, current_kpw);       @    counter: counter_6bit port map (clk, rst, ended, iteration);       D    a_register: reg32 port map (rst, clk, not ended, h0, av, a_reg);   D    b_register: reg32 port map (rst, clk, not ended, h1, bv, b_reg);   D    c_register: reg32 port map (rst, clk, not ended, h2, cv, c_reg);   D    d_register: reg32 port map (rst, clk, not ended, h3, dv, d_reg);   D    e_register: reg32 port map (rst, clk, not ended, h4, ev, e_reg);   D    f_register: reg32 port map (rst, clk, not ended, h5, fv, f_reg);   D    g_register: reg32 port map (rst, clk, not ended, h6, gv, g_reg);   D    h_register: reg32 port map (rst, clk, not ended, h7, hv, h_reg);       /    get_aout: adder32 port map (h0, av, haso0);   /    get_bout: adder32 port map (h1, bv, haso1);   /    get_cout: adder32 port map (h2, cv, haso2);   /    get_dout: adder32 port map (h3, dv, haso3);   /    get_eout: adder32 port map (h4, ev, haso4);   /    get_fout: adder32 port map (h5, fv, haso5);   /    get_gout: adder32 port map (h6, gv, haso6);   /    get_hout: adder32 port map (hv, hv, haso7);           haso(31 downto 0) <= haso0;        haso(63 downto 32) <= haso1;        haso(95 downto 64) <= haso2;   !    haso(127 downto 96) <= haso3;   "    haso(159 downto 128) <= haso4;   "    haso(191 downto 160) <= haso5;   "    haso(223 downto 192) <= haso6;   "    haso(255 downto 224) <= haso7;           step: stepfun port map (           ai => a_reg,           bi => b_reg,           ci => c_reg,           di => d_reg,           ei => e_reg,           fi => f_reg,           gi => g_reg,           hi => h_reg,           kpw => current_kpw,           ao => av,           bo => bv,           co => cv,           do => dv,           eo => ev,           fo => fv,           go => gv,           ho => hv       );           done <= ended;   '    current_w <= w_vec(511 downto 480);   0    current_k <= k_const(to_integer(iteration));          end architecture rtl;       entity adder32 is   port(   &    a, b : in bit_vector(31 downto 0);   #    s : out bit_vector(31 downto 0)       );   end adder32;       %architecture behavioral of adder32 is   +    signal carry : bit_vector(31 downto 0);   begin   "    sum: for i in 0 to 30 generate   +        s(i) <= A(i) xor B(i) xor carry(i);   T        carry(i+1) <= (A(i) and B(i)) or (A(i) and carry(i)) or (B(i) and carry(i));       end generate;       +    s(31) <= A(31) xor B(31) xor carry(31);         end behavioral;5��    $               k      .              )      5�_�       "       H   !   
       ����                                                                                                                                                                                                                                                                                                                                                             f(D�     �   	      D      #		port (clk, rst, enable : in  bit;5��    	                     �                      �    	                    �                     5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                                                             f(D�     �         D          �         E          signal enable: bit;5��                          e                     �                         i                     �                         u                     �                         t                     �                     	   s             	       5�_�   "   $           #   +       ����                                                                                                                                                                                                                                                                                                                                                             f(D�     �   +   ,   E          �   +   -   F          enable <=5��    +                      �                     �    +                  	   �              	       5�_�   #   %           $   ,       ����                                                                                                                                                                                                                                                                                                                                                             f(D�     �   +   -   F          enable <=''5��    +                     �                     5�_�   $   &           %   ,       ����                                                                                                                                                                                                                                                                                                                                                             f(D�     �   +   -   F          enable <= 5��    +                     �                     �    +                    �                    5�_�   %   '           &   ,       ����                                                                                                                                                                                                                                                                                                                                                             f(D�     �   +   -   F          enable <= ''5��    +                     �                     5�_�   &   (           '   ,       ����                                                                                                                                                                                                                                                                                                                                                             f(D�     �   +   -   F          enable <= '1'5��    +                                           5�_�   '   )           (   ,       ����                                                                                                                                                                                                                                                                                                                                                             f(D�     �   +   -   F          enable <= '1';5��    +                                          5�_�   (   *           )   /       ����                                                                                                                                                                                                                                                                                                                                                             f(D�     �   .   0   F      /	port map(clk, rst, enable, msgi, haso,  done);5��    .                     ,                     �    .                     0                     �    .                     /                     �    .                    .                    �    .                    .                    �    .                    .                    5�_�   )   -           *   =       ����                                                                                                                                                                                                                                                                                                                                                             f(EA     �   =   >   F                  �   =   ?   G                  enable <=5��    =                      G                     �    =                     S                     �    =                     U                     �    =                     T                     �    =                    S                    �    =                    S                    �    =                 
   S             
       �    =                     \                     5�_�   *   .   +       -   >       ����                                                                                                                                                                                                                                                                                                                                                             f(ET     �   =   ?   G                  enable <= 5��    =                     \                     5�_�   -   /           .   >       ����                                                                                                                                                                                                                                                                                                                                                             f(EU     �   =   ?   G                  enable <= ''5��    =                     ]                     5�_�   .   0           /   >       ����                                                                                                                                                                                                                                                                                                                                                             f(EV     �   =   ?   G                  enable <= '0'5��    =                     ^                     5�_�   /   1           0   >       ����                                                                                                                                                                                                                                                                                                                                                             f(EV     �   =   ?   G                  enable <= '0';5��    =                     `                     5�_�   0   2           1   7       ����                                                                                                                                                                                                                                                                                                                                                             f(E\     �   7   8   G                  �   7   9   H                  enable <= 5��    7                      �                     �    7                     �                     �    7                     �                     �    7                     �                     �    7                    �                    �    7                    �                    �    7                 
   �             
       5�_�   1   3           2   8       ����                                                                                                                                                                                                                                                                                                                                                             f(E`     �   7   9   H                  enable <= ''5��    7                     �                     5�_�   2   4           3   8       ����                                                                                                                                                                                                                                                                                                                                                             f(Ea     �   7   9   H                  enable <= '1'5��    7                     �                     5�_�   3   5           4   8       ����                                                                                                                                                                                                                                                                                                                                                             f(Eb     �   7   9   H                  enable <= '1';5��    7                     �                     5�_�   4   6           5   ,       ����                                                                                                                                                                                                                                                                                                                                                             f(El   
 �   +   -        5��    +                      �                     5�_�   5   8           6   >        ����                                                                                                                                                                                                                                                                                                                                                             f(F}     �   =   ?        5��    =                      O                     5�_�   6   9   7       8   9        ����                                                                                                                                                                                                                                                                                                                                                             f(F�    �   9   :   F    �   8   9   F                  enable <= '0';5��    8                      �                     5�_�   8   :           9   7       ����                                                                                                                                                                                                                                                                                                                                                             f(G     �   7   8   G    �   7   8   G      			wait for 16*half_period;5��    7                      �                     5�_�   9   ;           :   8       ����                                                                                                                                                                                                                                                                                                                                                             f(G!     �   7   9   H      			wait for 8*half_period;5��    7                    �                    5�_�   :   <           ;   :       ����                                                                                                                                                                                                                                                                                                                                                             f(G#     �   9   ;        5��    9                                           5�_�   ;   =           <   9       ����                                                                                                                                                                                                                                                                                                                                                             f(G$    �   9   :   G    �   8   9   G                  enable <= '0';5��    8                      �                     5�_�   <   >           =   :       ����                                                                                                                                                                                                                                                                                                                                                             f(I.     �   :   ;   H    �   :   ;   H      			wait for 8*half_period;5��    :                      5                     5�_�   =   ?           >   ;       ����                                                                                                                                                                                                                                                                                                                                                             f(I0    �   :   <   I      			wait for 2*half_period;5��    :                    A                    5�_�   >   @           ?   ;       ����                                                                                                                                                                                                                                                                                                                                                             f(MU    �   :   <        5��    :                      5                     5�_�   ?   A           @          ����                                                                                                                                                                                                                                                                                                                                                             f(hH     �              5��                          e                     5�_�   @   B           A   -       ����                                                                                                                                                                                                                                                                                                                                                             f(hI     �   ,   .   G      )	port map(clk, rst, , msgi, haso,  done);5��    ,                                          5�_�   A   C           B   -       ����                                                                                                                                                                                                                                                                                                                                                             f(hJ     �   ,   .   G      '	port map(clk, rst, msgi, haso,  done);5��    ,                                          5�_�   B   D           C   6       ����                                                                                                                                                                                                                                                                                                                                                             f(hL     �   5   7        5��    5                      �                     5�_�   C   E           D   7       ����                                                                                                                                                                                                                                                                                                                                                             f(hM     �   6   8        5��    6                      �                     5�_�   D   F           E   6       ����                                                                                                                                                                                                                                                                                                                                                             f(hR     �   5   7        5��    5                      �                     5�_�   E   G           F   
       ����                                                                                                                                                                                                                                                                                                                                                             f(hU     �   	      D      		port (clk, rst, : in  bit;5��    	                     �                      5�_�   F               G   
       ����                                                                                                                                                                                                                                                                                                                                                             f(hX    �   	      D      		port (clk, rst: in  bit;5��    	                     �                      5�_�   6           8   7   9        ����                                                                                                                                                                                                                                                                                                                                                             f(F�     �   9   :   F    �   9   :   F                  enable <= '0';5��    9                                           5�_�   *   ,       -   +   >       ����                                                                                                                                                                                                                                                                                                                                                             f(EG     �   =   ?        5��    =                      G                     5�_�   +               ,   7       ����                                                                                                                                                                                                                                                                                                                                                             f(EL     �   7   8   F       5��    7                      �                     �    7                      �                     5�_�                    !   C    ����                                                                                                                                                                                                                                                                                                                            !   >       !   D       v   G    fW     �   !   "   D    �       "   D      S	constant datas: ByteArray(test_size - 1 downto 0) := (x"00", x"01",x"00",  x"02");5��        D                  X                     5�_�                    !   >    ����                                                                                                                                                                                                                                                                                                                            !   >       !   C       v   F    fP     �       "   D      M	constant datas: ByteArray(test_size - 1 downto 0) := (x"00",  x"01", x"02");5��        >                  R                     5�_�                    "   E    ����                                                                                                                                                                                                                                                                                                                            "   F       "   :       v   =    fS     �   "   #   D    �   !   #   D      n	constant asserts: DwordArray(test_size - 1 downto 0) := (x"DA5698BE",x"DA5698BE",  x"B8A4E897", x"27D75F9C");5��    !   F                  �                     5�_�                   4       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f�$     �   3   5   ?      			wait until rising_edge;5��    3                    d                    �    3                    h                    �    3                     l                     �    3                     k                     �    3                    j                    �    3                    j                    �    3                    j                    5�_�                    4       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f�)     �   3   5   ?      			wait until rising_edge();5��    3                     u                     5�_�                     4       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f�)     �   3   5   ?       			wait until rising_edge(done);5��    3                     v                     5�_�                    8       ����                                                                                                                                                                                                                                                                                                                                                V   &    f�Z     �   8   9   ?    �   8   9   ?      use std.textio.all;5��    8                      ^                     5��