Vim�UnDo� V_KD�cx��ֽ]�xG�Ϛ[QZ�Mb~��_�   o           !                   e���    _�                           ����                                                                                                                                                                                                                                                                                                                                                             e��     �         �       �         �    �         �    5��                          (                      �                          (                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             e��    �                 5��                          E                      5�_�                    G       ����                                                                                                                                                                                                                                                                                                                                                             e���     �   F   H   �      P    signal convertedIn1: signed(32 downto 0); -- entrada convertida para 33 bits5��    F                     �                     5�_�                    G        ����                                                                                                                                                                                                                                                                                                                                                             e���     �   F   H   �      R    signal convertedIn1: signed()(32 downto 0); -- entrada convertida para 33 bits5��    F                      �                     5�_�                    G   +    ����                                                                                                                                                                                                                                                                                                                                                             e���     �   F   H   �      Q    signal convertedIn1: signed((32 downto 0); -- entrada convertida para 33 bits�   G   H   �    5��    F   ,                  �                     5�_�      	              G        ����                                                                                                                                                                                                                                                                                                                                                             e���     �   F   H   �      R    signal convertedIn1: signed((32 downto 0)); -- entrada convertida para 33 bits5��    F                      �                     �    F                     �                    �    F                  
   �             
       �    F           
       
   �      
       
       �    F           
          �      
              �    F                  
   �             
       5�_�                 	          ����                                                                                                                                                                                                                                                                                                                                                             e��}     �                use IEEE.std_logic_1164.ALL;5��                          (                      5�_�   	      
          $        ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �   $   (   �    �   $   %   �    5��    $                      �              )       5�_�                   3        ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �   3   7   �    �   3   4   �    5��    3                      �              )       5�_�                    B        ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �   B   F   �    �   B   C   �    5��    B                      �              )       5�_�                   O       ����                                                                                                                                                                                                                                                                                                                                                  V        e���     �   N   P   �      \    signal convertedIn1: signed(bit_vector(32 downto 0)); -- entrada convertida para 33 bits5��    N                     �                     5�_�                    O       ����                                                                                                                                                                                                                                                                                                                                                  V        e���     �   N   P   �      [    signal convertedIn1: signedbit_vector(32 downto 0)); -- entrada convertida para 33 bits5��    N          
           �      
               5�_�                    O   +    ����                                                                                                                                                                                                                                                                                                                                                  V        e���     �   N   P   �      Q    signal convertedIn1: signed(32 downto 0)); -- entrada convertida para 33 bits5��    N   +                  �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                       B           V        e��     �              B   library ieee;   use ieee.numeric_bit.all;       entity ch is   	port (   )    	x, y, z: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end ch;       architecture arch1 of ch is   0	signal op1, op2, op3 : bit_vector(31 downto 0);   begin   	op1 <= x and y;       op2 <= (not x) and z;       op3 <= op1 xor op2;        q <= op3;   
end arch1;       entity maj is   	port (   )    	x, y, z: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end maj;       architecture arch2 of maj is   4	signal op1, op2, op3, op4: bit_vector(31 downto 0);   begin   	op1 <= x and y;       op2 <= x and z;       op3 <= y and z;        op4 <= op1 xor op2 xor op3;        q <= op4;   
end arch2;       library ieee;   use ieee.numeric_bit.all;       entity sum0 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   	end sum0;       architecture arch3 of sum0 is   begin   1    q <= (x ror 2) xor (x ror 13) xor (x ror 22);   
end arch3;       library ieee;   use ieee.numeric_bit.all;       entity sum1 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   	end sum1;       architecture arch4 of sum1 is   begin   1    q <= (x ror 6) xor (x ror 11) xor (x ror 25);   
end arch4;    5��            B                       �              5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        e��r     �         [       �         [    �         Z    5��                          (                      �                         (               l       5�_�                       #    ����                                                                                                                                                                                                                                                                                                                                                  V        e��u     �         ^      #use IEEE.std_logic_unsigned.all; or5��       "                  u                      �                          s                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        e��z     �                use ieee.numeric_bit.all;5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        e��{     �         ]    �         ]    5��                                                5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        e��|     �                 library ieee;5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �         ]      use IEEE.std_logic_1164.all;    use IEEE.std_logic_unsigned.all;   use IEEE.std_logic_arith.all;5��                         (       \       e       5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �         ]      -- use IEEE.std_logic_1164.all;5��                         (                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �                use IEEE.std_logic_1164.all;5��                          (                      5�_�                             ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �         \      #-- use IEEE.std_logic_unsigned.all;5��                         (       $       !       5�_�      !                       ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �                 use IEEE.std_logic_unsigned.all;5��                          (       !               5�_�       "           !           ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �         [       -- use IEEE.std_logic_arith.all;5��                         (       !              5�_�   !   #           "           ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �                use IEEE.std_logic_arith.all;5��                          (                      5�_�   "   $           #           ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �         ^      use IEEE.numeric_std.all;�         \      ieee�         [       �         Z    5��                          (                      �                          (                      �                          )                      �                         +                      �                         *                      �                         )                     �                         )                     �                         )                     �                          )                      �                         )               D       �                          m                       5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �                use ieee.numeric_bit.all;5��                                                5�_�   $   &           %           ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �         ]    �         ]    5��                                                5�_�   %   '           &           ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �                 library IEEE;    5��                                                  5�_�   &   (           '           ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �         \      use ieee.numeric_bit.all;5��                                              5�_�   '   )           (           ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �         \      -- use ieee.numeric_bit.all;5��                                              5�_�   (   *           )           ����                                                                                                                                                                                                                                                                                                                                                  V        e���     �         \      use ieee.numeric_bit.all;5��                                              5�_�   )   +           *           ����                                                                                                                                                                                                                                                                                                                                                  V        e���     �         \      use IEEE.std_logic_1164.all;5��                         +                      5�_�   *   ,           +           ����                                                                                                                                                                                                                                                                                                                                                  V        e���     �         \      -- use IEEE.std_logic_1164.all;5��                         +                      5�_�   +   -           ,           ����                                                                                                                                                                                                                                                                                                                                                  V        e���     �         \      use IEEE.numeric_std.all;5��                         H                     5�_�   ,   .           -           ����                                                                                                                                                                                                                                                                                                                                                  V        e���     �         \      -- use IEEE.numeric_std.all;5��                         H                     5�_�   -   /           .           ����                                                                                                                                                                                                                                                                                                                                                  V        e���     �                use IEEE.numeric_std.all;5��                          H                      5�_�   .   0           /           ����                                                                                                                                                                                                                                                                                                                                                  V        e���     �         [      -- use ieee.numeric_bit.all;5��                                              5�_�   /   1           0           ����                                                                                                                                                                                                                                                                                                                                                  V        e���    �                use IEEE.std_logic_1164.all;5��                          (                      5�_�   0   2           1           ����                                                                                                                                                                                                                                                                                                                                                  V        e�S     �      
   Z    �      	   Z    5��                          �               D       5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                                                  V        e�T     �                C        a0, b0, c0, d0, e0, f0, g0, h0: out bit_vector(31 downto 0)5��                          �       D               5�_�   2   4           3   <        ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �   X   Z              h0 <= hi;�   W   Y              g0 <= gi;�   V   X              f0 <= fi;�   U   W              e0 <= preOut1(31 downto 0);�   T   V              d0 <= di;�   S   U              c0 <= ci;�   R   T              b0 <= bi;�   Q   S              a0 <= preOut2(31 downto 0);�   G   I          O    convertedIn5 <= signed('0' & ch01); -- extensão de sinal: número positivo�   ;   =   Z      $        port map (ei, fi, gi, ch01);5��    ;                    "                    �    G   "                 
                    �    Q                    �                    �    R                                        �    S                                        �    T                    '                    �    U                    5                    �    V                    U                    �    W                    c                    �    X                    q                    5�_�   3   5           4   "        ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �   !   "              component ch is           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;    5��    !                      �      �               5�_�   4   6           5           ����                                                                                                                                                                                                                                                                                                                                                  V        e�      �      "   S    �         S    5��                          /              �       5�_�   5   8           6   0        ����                                                                                                                                                                                                                                                                                                                                                  V        e�     �   /   0              component maj is           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;    5��    /                            �               5�_�   6   9   7       8   !        ����                                                                                                                                                                                                                                                                                                                                                  V        e�     �   !   )   S    �   !   "   S    5��    !                      �              �       5�_�   8   :           9   )        ����                                                                                                                                                                                                                                                                                                                                                  V        e�
     �   (   )              component sum1 is           port (   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;    5��    (                      l      �               5�_�   9   ;           :   /        ����                                                                                                                                                                                                                                                                                                                                                  V        e�     �   /   7   S    �   /   0   S    5��    /                                    �       5�_�   :   <           ;   Z       ����                                                                                                                                                                                                                                                                                                                                                  V        e�C     �   _              end entity �   [   ]   `      
entity  is�   ]                      �   [              ent�   Z               �   Z            5��    Z                      �                     �    Z                      �                     �    [                      �                     �    [                    �                    �    [                     �                     �    [                     �                     �    [                     �                     �    [                     �                     �    [                     �                    �    [                     �                     �    [                     �                     �    [                     �                    �    [                     �                    �    [                     �                    �    [                     �                    �    [                    �                     �    ]                      �                      �    ]                    �                     �    _                     �                     �    [                     �                     �    _                     �                     5�_�   ;   =           <   \       ����                                                                                                                                                                                                                                                                                                                            \   
       \          v       e�K     �   ]   _   `              �   \   ]   `    �   _              end entity exp3;�   [   ]   `      entity exp3 is�   \   ]   `    �   \   ]   `    �   \   ]   `    �   \   ]   `    5��    [                    �                    �    _                    �                    �    [                     �                     �    _                    �                    �    [   	                  �                     �    _                    �                    �    [   
                  �                     �    _                    �                    �    [   
                  �                     �    [   	                  �                     �    [                     �                     �    [                    �                    �    [                    �                    �    [                    �                    �    _                    �                    �    ]                     �                     �    ]                 	   �             	       �    ]                     �                     �    ]                     �                     �    ]                 
   �             
       �    ]          
          �      
              �    ]                 
   �             
       5�_�   <   >           =   ^       ����                                                                                                                                                                                                                                                                                                                            \   
       \          v       e�[     �   ]   _   `              A: in bit_vector5��    ]                     �                     5�_�   =   ?           >   ^       ����                                                                                                                                                                                                                                                                                                                            \   
       \          v       e�]     �   ]   _   `              A: in bit_vector()5��    ]                     �                     �    ]                    �                    �    ]                    �                    �    ]                    �                    5�_�   >   @           ?   ^   %    ����                                                                                                                                                                                                                                                                                                                            \   
       \          v       e�a     �   ]   _   `      %        A: in bit_vector(31 downto 0)5��    ]   %                  �                     �    ]   %                 �                    �    ]   %                 �                    �    ]   %                 �                    5�_�   ?   B           @   ^   %    ����                                                                                                                                                                                                                                                                                                                            \   
       \          v       e�f     �   ^   `   `    �   ^   _   `    5��    ^                      �              '       5�_�   @   C   A       B   _   %    ����                                                                                                                                                                                                                                                                                                                            \   
       \          v       e�i     �   _   a   a    �   _   `   a    5��    _                      �              '       5�_�   B   D           C   `       ����                                                                                                                                                                                                                                                                                                                            \   
       \          v       e�k     �   _   a   b      &        A: in bit_vector(31 downto 0);5��    _                    �                    5�_�   C   E           D   _       ����                                                                                                                                                                                                                                                                                                                            \   
       \          v       e�l     �   ^   `   b      &        A: in bit_vector(31 downto 0);5��    ^                    �                    5�_�   D   F           E   `   %    ����                                                                                                                                                                                                                                                                                                                            \   
       \          v       e�n     �   _   a   b      &        S: in bit_vector(31 downto 0);5��    _   %                                       5�_�   E   G           F   ^   	    ����                                                                                                                                                                                                                                                                                                                            `          ^                 e�}     �   ^   a   b      &        B: in bit_vector(31 downto 0);   %        S: in bit_vector(31 downto 0)�   ]   _   b      &        A: in bit_vector(31 downto 0);5��    ]   	                  �                     �    ^   	                  �                     �    _   	                  �                     5�_�   F   H           G   `       ����                                                                                                                                                                                                                                                                                                                            `          ^                 e��     �   _   a   b      &        S : in bit_vector(31 downto 0)5��    _                                         5�_�   G   I           H   b       ����                                                                                                                                                                                                                                                                                                                            `          ^                 e��     �   i              end architecture �   c   e   j      architecture rtl of  is�   g                  �   c              arch�   b               �   b            5��    b                      7                     �    b                      7                     �    c                      8                     �    c                     ;                     �    c                     :                     �    c                     9                     �    c                     8                    �    c                     8                    �    c                     8                    �    c                     8                    �    c                    L                     �    g                      d                      �    g                    d                     �    i                     {                     �    c                     L                     �    i                                          5�_�   H   J           I   e        ����                                                                                                                                                                                                                                                                                                                            d          j          V       e��     �   i              end architecture �   c   e   j      architecture rtl of  is�   g                  �   c              architecture rtl of exp3 is�   d   e                 begin                        end architecture rtl;5��    d                      T      0               �    c                     8                    �    c                     ;                     �    c                     :                     �    c                     9                     �    c                     8                    �    c                     8                    �    c                     8                    �    c                     8                    �    c                    L                     �    g                      d                      �    g                    d                     �    i                     {                     �    c                     L                     �    i                                          5�_�   I   K           J   d       ����                                                                                                                                                                                                                                                                                                                            d          d          v       e��     �   d   e   j    �   i              end architecture rtl;�   d   e   j    �   d   e   j    �   d   e   j    �   d   e   j    �   d   e   j    �   d   e   j    �   d   e   j    �   d   e   j    �   d   e   j    �   c   e   j      architecture rtl of exp3 is5��    c                    E                    �    i                    }                    �    c                     F                     �    i                    ~                    �    c                     G                     �    i                                        �    c                     H                     �    i                    �                    �    c                     I                     �    i                    �                    �    c                     J                     �    i                    �                    �    c                     K                     �    i                    �                    �    c                     L                     �    i                    �                    �    c                     M                     �    i                 	   �             	       �    c                     N                     �    i          	       
   �      	       
       5�_�   J   L           K   d       ����                                                                                                                                                                                                                                                                                                                            d          d          v       e��     �   g   i   j          �   c   e   j      "architecture behavioral of exp3 is5��    c                    S                    �    c                     U                     �    c                     T                     �    c                    S                    �    c                    S                    �    c                    S                    �    g                     r                     5�_�   K   M           L   h       ����                                                                                                                                                                                                                                                                                                                            d          d          v       e� �     �   h   s   j    �   h   i   j    5��    h               
       v              �      5�_�   L   N           M   g       ����                                                                                                                                                                                                                                                                                                                            d          d          v       e� �     �   f   g                     dwa5��    f                      i                     5�_�   M   O           N   e       ����                                                                                                                                                                                                                                                                                                                            d          d          v       e� �     �   d   e                 begin5��    d                      ^                     5�_�   N   P           O   h       ����                                                                                                                                                                                                                                                                                                                            d          d          v       e� �     �   g   i   p      &    gen_sum: for i in 0 to 30 generate5��    g                     �                     5�_�   O   S           P   h       ����                                                                                                                                                                                                                                                                                                                            d          d          v       e� �     �   g   i   p          : for i in 0 to 30 generate5��    g                     �                     5�_�   P   T   R       S   g       ����                                                                                                                                                                                                                                                                                                                            d          d          v       e�!     �   f   h   p      1    carry(0) <= '0';  -- inicialização do carry5��    f                     �                     5�_�   S   U           T   i   +    ����                                                                                                                                                                                                                                                                                                                            d          d          v       e�!     �   h   j   p      H        S(i) <= A(i) xor B(i) xor carry(i);  -- somando bits individuais5��    h   +                  �                     5�_�   T   V           U   j   T    ����                                                                                                                                                                                                                                                                                                                            d          d          v       e�!     �   i   k   p      j        carry(i+1) <= (A(i) and B(i)) or (A(i) and carry(i)) or (B(i) and carry(i));  -- atualizando carry5��    i   T                  C                     5�_�   U   W           V   m   ,    ����                                                                                                                                                                                                                                                                                                                            d          d          v       e�!     �   l   m          -    -- último bit soma sem atualizar o carry5��    l                      W      .               5�_�   V   X           W   Z        ����                                                                                                                                                                                                                                                                                                                                       Z           V        e�(6    �      [   o   W   entity stepfun is   
    port (   @    	ai, bi, ci, di, ei, fi, gi, hi: in bit_vector(31 downto 0);   (        kpw: in bit_vector(31 downto 0);   C        ao, bo, co, do, eo, fo, go, ho: out bit_vector(31 downto 0)   
        );   end stepfun;        architecture arch7 of stepfun is   P    signal convertedIn1: signed(32 downto 0); -- entrada convertida para 33 bits   P    signal convertedIn2: signed(32 downto 0); -- entrada convertida para 33 bits   P    signal convertedIn3: signed(32 downto 0); -- entrada convertida para 33 bits   P    signal convertedIn4: signed(32 downto 0); -- entrada convertida para 33 bits   P    signal convertedIn5: signed(32 downto 0); -- entrada convertida para 33 bits   P    signal convertedIn6: signed(32 downto 0); -- entrada convertida para 33 bits   P    signal convertedIn7: signed(32 downto 0); -- entrada convertida para 33 bits   P    signal convertedIn8: signed(32 downto 0); -- entrada convertida para 33 bits   J    signal internal1: signed(32 downto 0);     -- somador interno: 33 bits   J    signal internal2: signed(32 downto 0);     -- somador interno: 33 bits   `    signal preOut1: bit_vector(32 downto 0);  -- pré-saida: internal convertido para bit_vector   `    signal preOut2: bit_vector(32 downto 0);  -- pré-saida: internal convertido para bit_vector       -- Declaração dos componentes       component ch is           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component maj is           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component sum0 is           port (   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component sum1 is           port (   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;       begin       -- Saida dos Componentes       first: sum1           port map (ei, sum1_01);       second: ch    $        port map (ei, fi, gi, cho1);       third: sum0            port map (ai, sum0_01);       fourty: maj    $        port map (ai, bi, ci, maj1);           -- Somadores       M    convertedIn1 <= signed('0' & di); -- extensão de sinal: número positivo   M    convertedIn2 <= signed('0' & hi); -- extensão de sinal: número positivo   N    convertedIn3 <= signed('0' & kpw); -- extensão de sinal: número positivo   R    convertedIn4 <= signed('0' & sum1_01); -- extensão de sinal: número positivo   O    convertedIn5 <= signed('0' & cho1); -- extensão de sinal: número positivo   R    convertedIn6 <= signed('0' & sum0_01); -- extensão de sinal: número positivo   O    convertedIn7 <= signed('0' & maj1); -- extensão de sinal: número positivo       Z    internal1 <= convertedIn1 + convertedIn2 + convertedIn3 + convertedIn4 + convertedIn5;   i    internal2 <= convertedIn2 + convertedIn3 + convertedIn4 + convertedIn5 + convertedIn6 + convertedIn7;       %    preOut1 <= bit_vector(internal1);   %    preOut2 <= bit_vector(internal2);           ao <= preOut2(31 downto 0);       bo <= bi;       co <= ci;       do <= di;       eo <= preOut1(31 downto 0);       fo <= fi;       go <= gi;       ho <= hi;   
end arch7;5��           W       W       )       ]      W      5�_�   W   Y           X   h       ����                                                                                                                                                                                                                                                                                                                                       Z           V        e�(I    �   g   i   o          for i in 0 to 30 generate5��    g                     �                     5�_�   X   Z           Y          ����                                                                                                                                                                                                                                                                                                                            Z                    V       e�(Z    �      [   o   W   -- entity stepfun is   --     port (   C--     	ai, bi, ci, di, ei, fi, gi, hi: in bit_vector(31 downto 0);   +--         kpw: in bit_vector(31 downto 0);   F--         ao, bo, co, do, eo, fo, go, ho: out bit_vector(31 downto 0)   --         );   -- end stepfun;   --   #-- architecture arch7 of stepfun is   S--     signal convertedIn1: signed(32 downto 0); -- entrada convertida para 33 bits   S--     signal convertedIn2: signed(32 downto 0); -- entrada convertida para 33 bits   S--     signal convertedIn3: signed(32 downto 0); -- entrada convertida para 33 bits   S--     signal convertedIn4: signed(32 downto 0); -- entrada convertida para 33 bits   S--     signal convertedIn5: signed(32 downto 0); -- entrada convertida para 33 bits   S--     signal convertedIn6: signed(32 downto 0); -- entrada convertida para 33 bits   S--     signal convertedIn7: signed(32 downto 0); -- entrada convertida para 33 bits   S--     signal convertedIn8: signed(32 downto 0); -- entrada convertida para 33 bits   M--     signal internal1: signed(32 downto 0);     -- somador interno: 33 bits   M--     signal internal2: signed(32 downto 0);     -- somador interno: 33 bits   c--     signal preOut1: bit_vector(32 downto 0);  -- pré-saida: internal convertido para bit_vector   c--     signal preOut2: bit_vector(32 downto 0);  -- pré-saida: internal convertido para bit_vector   --   "-- -- Declaração dos componentes   --     component ch is   --         port (   3--             x, y, z: in bit_vector(31 downto 0);   ---             q: out bit_vector(31 downto 0)   --         );   --     end component;   --   --     component maj is   --         port (   3--             x, y, z: in bit_vector(31 downto 0);   ---             q: out bit_vector(31 downto 0)   --         );   --     end component;   --   --     component sum0 is   --         port (   ---             x: in bit_vector(31 downto 0);   ---             q: out bit_vector(31 downto 0)   --         );   --     end component;   --   --     component sum1 is   --         port (   ---             x: in bit_vector(31 downto 0);   ---             q: out bit_vector(31 downto 0)   --         );   --     end component;   --   -- begin   --     -- Saida dos Componentes   --     first: sum1   "--         port map (ei, sum1_01);   --     second: ch    '--         port map (ei, fi, gi, cho1);   --     third: sum0    "--         port map (ai, sum0_01);   --     fourty: maj    '--         port map (ai, bi, ci, maj1);   --   --     -- Somadores   --   P--     convertedIn1 <= signed('0' & di); -- extensão de sinal: número positivo   P--     convertedIn2 <= signed('0' & hi); -- extensão de sinal: número positivo   Q--     convertedIn3 <= signed('0' & kpw); -- extensão de sinal: número positivo   U--     convertedIn4 <= signed('0' & sum1_01); -- extensão de sinal: número positivo   R--     convertedIn5 <= signed('0' & cho1); -- extensão de sinal: número positivo   U--     convertedIn6 <= signed('0' & sum0_01); -- extensão de sinal: número positivo   R--     convertedIn7 <= signed('0' & maj1); -- extensão de sinal: número positivo   --   ]--     internal1 <= convertedIn1 + convertedIn2 + convertedIn3 + convertedIn4 + convertedIn5;   l--     internal2 <= convertedIn2 + convertedIn3 + convertedIn4 + convertedIn5 + convertedIn6 + convertedIn7;   --   (--     preOut1 <= bit_vector(internal1);   (--     preOut2 <= bit_vector(internal2);   --   "--     ao <= preOut2(31 downto 0);   --     bo <= bi;   --     co <= ci;   --     do <= di;   "--     eo <= preOut1(31 downto 0);   --     fo <= fi;   --     go <= gi;   --     ho <= hi;   -- end arch7;5��           W       W       )       W      ]      5�_�   Y   [           Z   ?       ����                                                                                                                                                                                                                                                                                                                            Z                    V       e��     �   >   @   o          fourty: maj 5��    >                    a                    5�_�   Z   \           [   S   
    ����                                                                                                                                                                                                                                                                                                                            Z                    V       e��B     �   R   T   o          bo <= bi;5��    R   
                                     5�_�   [   ]           \   T   
    ����                                                                                                                                                                                                                                                                                                                            Z                    V       e��K     �   S   U   o          co <= ci;5��    S   
                                     5�_�   \   ^           ]   U   
    ����                                                                                                                                                                                                                                                                                                                            Z                    V       e��Q     �   T   V   o          do <= di;5��    T   
                 -                    5�_�   ]   _           ^   W   
    ����                                                                                                                                                                                                                                                                                                                            Z                    V       e��X     �   V   X   o          fo <= fi;5��    V   
                 [                    5�_�   ^   `           _   X   
    ����                                                                                                                                                                                                                                                                                                                            Z                    V       e��_     �   W   Y   o          go <= gi;5��    W   
                 i                    5�_�   _   a           `   Y   
    ����                                                                                                                                                                                                                                                                                                                            Z                    V       e��d     �   X   Z   o          ho <= hi;5��    X   
                 w                    5�_�   `   b           a   5   
    ����                                                                                                                                                                                                                                                                                                                            Z                    V       e���     �   6   9   q          component�   5   8   p          �   5   7   o    5��    5                      �                     �    5                      �                     �    5                     �                     �    6                     �                     �    6                     �                     �    6                     �                     �    6                     �                     �    6                 	   �             	       �    6          	          �      	              �    6                    �                    �    6                    �                     �    7                     �                    5�_�   a   c           b   8       ����                                                                                                                                                                                                                                                                                                                            ]                    V       e���     �   7   9   r              port 5��    7                     �                     5�_�   b   d           c   8       ����                                                                                                                                                                                                                                                                                                                            ]                    V       e���     �   7   :   s              port (�   8   :                       )�   7   :   r              port ()5��    7                    �              	       �    8                     �                    �    7                    �              	       �    8                     �                     �    8                    �                    �    8                    �                    5�_�   c   e           d   9       ����                                                                                                                                                                                                                                                                                                                            e          c          V       e���     �   9   =   t    �   9   :   t    5��    9                      �              x       5�_�   d   f           e   9       ����                                                                                                                                                                                                                                                                                                                            h          f          V       e���     �   8   9                      A: in bi5��    8                      �                     5�_�   e   g           f   9       ����                                                                                                                                                                                                                                                                                                                            9          ;                 e���     �   9   <   v      '        B : in bit_vector(31 downto 0);   '        S : out bit_vector(31 downto 0)�   8   :   v      '        A : in bit_vector(31 downto 0);5��    8                     �                     �    9                     �                     �    :                     (                     5�_�   f   h           g   <       ����                                                                                                                                                                                                                                                                                                                            9          ;                 e���     �   ;   =   v                   )5��    ;                     X                     5�_�   g   i           h   <       ����                                                                                                                                                                                                                                                                                                                            9          ;                 e���     �   ;   =   v                  )5��    ;                     T                     5�_�   h   j           i   <   	    ����                                                                                                                                                                                                                                                                                                                            9          ;                 e���     �   <   >   w          end component�   ;   >   v      	        )5��    ;   	                  U                     �    ;   
                 V              	       �    <                     _                     �    <                     W                    �    <                     _                     �    <                     b                     �    <   
                  a                     �    <   	                  `                     �    <                 	   _             	       �    <          	          _      	              �    <                 
   _             
       5�_�   i   k           j   H       ����                                                                                                                                                                                                                                                                                                                            9          ;                 e���     �   H   K   x              �   H   J   w    5��    H                      Z	              	       �    H                      Z	                     �    H                     Z	              	       �    I                     c	                     �    I                    _	                    �    I                     `	                     �    I                    _	                    �    I                     `	                     �    I                     _	                     5�_�   j   l           k   B       ����                                                                                                                                                                                                                                                                                                                            9          ;                 e��(     �   @   B   y          first: sum1   port map (ei, sum1_01);�   A   C   y              port map (ei, sum1_01);5��    A                      �                     �    @                     �                     �    @                     �                     5�_�   k   m           l   C       ����                                                                                                                                                                                                                                                                                                                            9          ;                 e��,     �   A   C   x          second: ch    port map (ei, fi, gi, cho1);�   B   D   x      $        port map (ei, fi, gi, cho1);5��    B                      �                     �    A                     �                     5�_�   l   n           m   D       ����                                                                                                                                                                                                                                                                                                                            9          ;                 e��/     �   B   D   w          third: sum0    port map (ai, sum0_01);�   C   E   w              port map (ai, sum0_01);5��    C                      �                     �    B                     �                     5�_�   m   o           n   E       ����                                                                                                                                                                                                                                                                                                                            9          ;                 e��1     �   C   E   v          fourth: maj    port map (ai, bi, ci, maj1);�   D   F   v      $        port map (ai, bi, ci, maj1);5��    D                      	                     �    C                     	                     5�_�   n   p           o   E        ����                                                                                                                                                                                                                                                                                                                            9          ;                 e��4     �   E   G   u    �   E   F   u    5��    E                      8	              -       5�_�   o   q           p   G       ����                                                                                                                                                                                                                                                                                                                            9          ;                 e��6     �   F   G              5��    F                      e	                     5�_�   p   r           q   F       ����                                                                                                                                                                                                                                                                                                                            9          ;                 e��C     �   E   G   u      ,    fourth: maj port map (ai, bi, ci, maj1);5��    E                    <	                    5�_�   q   s           r   F       ����                                                                                                                                                                                                                                                                                                                            9          ;                 e��K     �   E   G   u      +    get_e: maj port map (ai, bi, ci, maj1);5��    E                     ?	                     5�_�   r   t           s   F       ����                                                                                                                                                                                                                                                                                                                            9          ;                 e��M     �   E   G   u      *    gete: maj port map (ai, bi, ci, maj1);5��    E                    ?	                    5�_�   s   u           t   F   
    ����                                                                                                                                                                                                                                                                                                                            9          ;                 e��N     �   E   G   u      *    getE: maj port map (ai, bi, ci, maj1);5��    E   
                 B	                    5�_�   t   v           u   F       ����                                                                                                                                                                                                                                                                                                                            9          ;                 e��[     �   E   G   u      .    getE: somador port map (ai, bi, ci, maj1);5��    E                    T	                    �    E                    U	                    �    E   "                  Z	                     �    E   !                 Y	                    �    E   %                 ]	                    �    E   %                 ]	                    �    E   %                 ]	                    5�_�   u   w           v      )    ����                                                                                                                                                                                                                                                                                                                            9          ;                 e���     �         u    �         u    5��                          �              Q       5�_�   v   x           w          ����                                                                                                                                                                                                                                                                                                                            :          <                 e���     �         v      P    signal convertedIn8: signed(32 downto 0); -- entrada convertida para 33 bits5��                        �                    5�_�   w   y           x          ����                                                                                                                                                                                                                                                                                                                            :          <                 e���     �         v    �         v    5��                                         J       5�_�   x   {           y          ����                                                                                                                                                                                                                                                                                                                            ;          =                 e���     �         w      I    signal chOut: signed(32 downto 0); -- entrada convertida para 33 bits5��                                            5�_�   y   |   z       {          ����                                                                                                                                                                                                                                                                                                                            ;          =                 e���     �         w    �         w    5��                          K              K       5�_�   {   }           |          ����                                                                                                                                                                                                                                                                                                                            <          >                 e���     �         x      J    signal majOut: signed(32 downto 0); -- entrada convertida para 33 bits5��                        V                    5�_�   |   ~           }          ����                                                                                                                                                                                                                                                                                                                            <          >                 e���     �         x    �         x    5��                          �              L       5�_�   }              ~          ����                                                                                                                                                                                                                                                                                                                            =          ?                 e���     �         y      K    signal sum0Out: signed(32 downto 0); -- entrada convertida para 33 bits5��                        �                    5�_�   ~   �                      ����                                                                                                                                                                                                                                                                                                                                                V       e���    �                K    signal sum1Out: signed(32 downto 0); -- entrada convertida para 33 bits�                K    signal sum0Out: signed(32 downto 0); -- entrada convertida para 33 bits�                J    signal majOut: signed(32 downto 0); -- entrada convertida para 33 bits�         y      I    signal chOut: signed(32 downto 0); -- entrada convertida para 33 bits5��                        �                    �                                            �                        g                    �                        �                    5�_�      �           �      '    ����                                                                                                                                                                                                                                                                                                                                                V       e���     �         y      I    signal chOut: signed(31 downto 0); -- entrada convertida para 33 bits5��       '       "           �      "               5�_�   �   �           �      (    ����                                                                                                                                                                                                                                                                                                                                                V       e���     �         y      J    signal majOut: signed(31 downto 0); -- entrada convertida para 33 bits5��       (       "                 "               5�_�   �   �           �      )    ����                                                                                                                                                                                                                                                                                                                                                V       e���     �         y      K    signal sum0Out: signed(31 downto 0); -- entrada convertida para 33 bits5��       )       "           0      "               5�_�   �   �           �      )    ����                                                                                                                                                                                                                                                                                                                                                V       e���     �         y      K    signal sum1Out: signed(31 downto 0); -- entrada convertida para 33 bits5��       )       "           Z      "               5�_�   �   �           �      &    ����                                                                                                                                                                                                                                                                                                                                                V       e���     �         z          �         y    5��                          �                     �                          �                     �                         �                     �                         �                     �       
                 �                    5�_�   �   �           �      !    ����                                                                                                                                                                                                                                                                                                                                                V       e���     �         {    5��                                               �                                               5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                                                V       e���     �   H   I          +    second: ch port map (ei, fi, gi, cho1);5��    H                      �	      ,               5�_�   �   �           �   H       ����                                                                                                                                                                                                                                                                                                                                                V       e���     �   G   I   {    �   H   I   {    5��    G                      X	              ,       5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                                                V       e���     �   J   K          ,    fourth: maj port map (ai, bi, ci, maj1);5��    J                      �	      -               5�_�   �   �           �   I        ����                                                                                                                                                                                                                                                                                                                                                V       e���     �   H   J   {    �   I   J   {    5��    H                      �	              -       5�_�   �   �           �   J       ����                                                                                                                                                                                                                                                                                                                                                V       e���     �   I   K   |      '    first: sum1 port map (ei, sum1_01);5��    I                     �	                     5�_�   �   �           �   H       ����                                                                                                                                                                                                                                                                                                                            H          H   	       v   	    e��     �   G   I   |      +    second: ch port map (ei, fi, gi, cho1);�   H   I   |    5��    G                    \	                    5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            I          I   	       v   	    e��     �   H   J   |      ,    fourth: maj port map (ai, bi, ci, maj1);�   I   J   |    5��    H                    �	                    5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                            K          K          v       e��     �   J   L   |      '    third: sum0 port map (ai, sum0_01);�   K   L   |    5��    J                    �	                    5�_�   �   �           �   J       ����                                                                                                                                                                                                                                                                                                                            K          K   	       v       e��     �   I   K   |      "    : sum1 port map (ei, sum1_01);�   J   K   |    5��    I                     �	                     5�_�   �   �           �   J       ����                                                                                                                                                                                                                                                                                                                            K          K   	       v       e��     �   I   J          '    third: sum1 port map (ei, sum1_01);5��    I                      �	      (               5�_�   �   �   �       �   J       ����                                                                                                                                                                                                                                                                                                                            J          J   	       v       e��     �   I   K   {    �   J   K   {    5��    I                      �	              (       5�_�   �   �           �   H   $    ����                                                                                                                                                                                                                                                                                                                            K          K   	       v       e��     �   G   I   |      *    first: ch port map (ei, fi, gi, cho1);5��    G   $                 |	                    �    G   %                  }	                     �    G   $                 |	                    �    G   '                  	                     �    G   &                  ~	                     �    G   %                  }	                     �    G   $                 |	                    �    G   (                  �	                     �    G   '                  	                     �    G   &                  ~	                     �    G   %                  }	                     �    G   $                 |	                    �    G   $                 |	                    �    G   $                 |	                    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��6     �                )    signal sum1Out: signed(31 downto 0); �                )    signal sum0Out: signed(31 downto 0); �                (    signal majOut: signed(31 downto 0); �         |      '    signal chOut: signed(31 downto 0); 5��                     
   �             
       �                     
                
       �                     
   G             
       �                     
   u             
       5�_�   �   �           �   I   &    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��=     �   H   J   |      ,    second: maj port map (ai, bi, ci, maj1);5��    H   &                 �	                    �    H   )                  �	                     �    H   (                  �	                     �    H   '                  �	                     �    H   &                 �	                    �    H   &                 �	                    �    H   &                 �	                    5�_�   �   �           �   J       ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��A     �   I   K   |      '    third: sum1 port map (ei, sum1_01);5��    I                    �	                    �    I                    �	                    �    I   !                  �	                     �    I                      �	                     �    I                     �	                     �    I                    �	                    �    I                    �	                    �    I                    �	                    5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��G     �   J   L   |      (    fourth: sum0 port map (ai, sum0_01);5��    J                    

                    �    J   #                  
                     �    J   "                  
                     �    J   !                  
                     �    J                      
                     �    J                    

                    �    J                    

                    �    J                    

                    5�_�   �   �           �   M   *    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �   L   N   |      ,    getE: somador port map (A => ei, B => );5��    L   *                  ?
                     �    L   -                  B
                     �    L   ,                  A
                     �    L   +                  @
                     �    L   *                 ?
                    �    L   -                  B
                     �    L   ,                  A
                     �    L   +                  @
                     �    L   *                 ?
                    �    L   *                 ?
                    �    L   *                 ?
                    �    L   *                 ?
                    5�_�   �   �           �   M   1    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �   L   N   |      3    getE: somador port map (A => ei, B => sum1Out);5��    L   1               	   F
              	       �    L   9                  N
                     �    L   8                 M
                    �    L   8                 M
                    �    L   8                 M
                    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �         |      `    signal preOut1: bit_vector(32 downto 0);  -- pré-saida: internal convertido para bit_vector5��                         F                    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �          |      `    signal preOut2: bit_vector(32 downto 0);  -- pré-saida: internal convertido para bit_vector5��                         �                    5�_�   �   �           �      ;    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �         |      `    signal preOut1: bit_vector(31 downto 0);  -- pré-saida: internal convertido para bit_vector5��       ;       %           a      %               5�_�   �   �           �      ;    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �         |      ;    signal preOut1: bit_vector(31 downto 0);  -- pré-saida5��       ;                  a                     5�_�   �   �           �      =    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �         |      =    signal preOut1: bit_vector(31 downto 0);  -- pré-saida e5��       =                  c                     5�_�   �   �           �      ;    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �          |      `    signal preOut2: bit_vector(31 downto 0);  -- pré-saida: internal convertido para bit_vector5��       ;       %           �      %               5�_�   �   �           �      ;    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �          |      ;    signal preOut2: bit_vector(31 downto 0);  -- pré-saida5��       ;                  �                     5�_�   �   �           �      <    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �         |      >    signal preOut1: bit_vector(31 downto 0);  -- pré-saida eo5��       <                 b                    5�_�   �   �           �      <    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �          |      >    signal preOut2: bit_vector(31 downto 0);  -- pré-saida ao5��       <                 �                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �         |      >    signal preOut1: bit_vector(31 downto 0);  -- pré-saida ao5��                        7                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �         |      A    signal preOutAout: bit_vector(31 downto 0);  -- pré-saida ao5��                         4                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �         |      >    signal preAout: bit_vector(31 downto 0);  -- pré-saida ao5��                        5                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �          |      >    signal preOut2: bit_vector(31 downto 0);  -- pré-saida eo5��                        s                    5�_�   �   �           �   M   8    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �   L   N   |      A    getE: somador port map (A => ei, B => sum1Out, S => preOut1);5��    L   8                 	
                    �    L   ;                 
                    �    L   ;                  
                     �    L   :                  
                     �    L   9                  

                     �    L   8                 	
                    �    L   8                 	
                    �    L   8                 	
                    5�_�   �   �           �   c   
    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �   b   d   |          eo <= preOut1(31 downto 0);5��    b   
                 �                    �    b                     �                     �    b                     �                     �    b                     �                     �    b   
                 �                    �    b   
                 �                    �    b   
                 �                    5�_�   �   �           �   c       ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �   b   d   |          eo <= preEOut(31 downto 0);5��    b                     �                     5�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��     �   M   O   |    �   M   N   |    5��    M                      
              B       5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��     �   M   O   }      A    getE: somador port map (A => ei, B => sum1Out, S => preEOut);5��    M                    
                    5�_�   �   �           �   N   $    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��     �   M   O   }      D    getChIn: somador port map (A => ei, B => sum1Out, S => preEOut);5��    M   $                 7
                    5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��0     �   M   O   }      D    getChIn: somador port map (A => hi, B => sum1Out, S => preEOut);5��    M                    
                    5�_�   �   �           �   N   2    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��B     �   M   O   }      I    chComplement: somador port map (A => hi, B => sum1Out, S => preEOut);5��    M   2                 E
                    5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��O     �   M   O   }      E    chComplement: somador port map (A => hi, B => kpw, S => preEOut);5��    M                     
                     �    M                    
                    5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��Q     �   M   O   }      H    getchComplement: somador port map (A => hi, B => kpw, S => preEOut);5��    M                    
                    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��_     �         ~          �         }    5��                          �                     �                          �                     �                          �                     �                         �                     �                          �                     5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��`     �             �             5��                          �              Q       5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��b     �         �       5��                          �                     �                          �                     5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��c     �         �       5��                          �                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��l     �         �      P    signal convertedIn8: signed(32 downto 0); -- entrada convertida para 33 bits5��                        �                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��s     �         �      P    signal chComplement: signed(32 downto 0); -- entrada convertida para 33 bits5��                        �                    �                         �                     �                         �                     �                     
   �             
       �              
          �      
              �                     
   �             
       5�_�   �   �           �      %    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��v     �         �      T    signal chComplement: bit_vector(32 downto 0); -- entrada convertida para 33 bits5��       %                 �                    5�_�   �   �           �      2    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��y     �         �      T    signal chComplement: bit_vector(31 downto 0); -- entrada convertida para 33 bits5��       2       "                 "               5�_�   �   �           �      1    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e��z     �         �      2    signal chComplement: bit_vector(31 downto 0); 5��       1                                        5�_�   �   �           �      0    ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �         �    �         �    5��                                        2       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �         �    �         �    5��                          3              2       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               &          (       V   (    e���     �         �    �         �    5��                          e              2       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       e���     �         �      1    signal chComplement: bit_vector(31 downto 0);5��                                            5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       e���     �                1    signal chComplement: bit_vector(31 downto 0);5��                          5      2               5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       e���     �         �    �         �    5��                                        2       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       e���     �         �      1    signal chComplement: bit_vector(31 downto 0);5��                                            5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       e���     �         �      1    signal chComplement: bit_vector(31 downto 0);5��                        s                    5�_�   �   �           �   T   ?    ����                                                                                                                                                                                                                                                                                                                                                v       e���     �   S   U   �      H    getChComplement: somador port map (A => hi, B => kpw, S => preEOut);5��    S   ?                 8                    �    S   A                  :                     �    S   @                  9                     �    S   ?                 8                    �    S   ?                 8                    �    S   ?                 8                    5�_�   �   �           �   T   J    ����                                                                                                                                                                                                                                                                                                                                                v       e���     �   T   V   �    �   T   U   �    5��    T                      G              N       5�_�   �   �           �   U       ����                                                                                                                                                                                                                                                                                                                            U          U          v       e���     �   T   V   �      M    getChComplement: somador port map (A => hi, B => kpw, S => chComplement);5��    T                    N                    5�_�   �   �           �   U   .    ����                                                                                                                                                                                                                                                                                                                            U          U          v       e���     �   T   V   �      O    getSum1Complement: somador port map (A => hi, B => kpw, S => chComplement);5��    T   .                 u                    �    T   1                  x                     �    T   0                  w                     �    T   /                  v                     �    T   .                 u                    �    T   .                 u                    �    T   .                 u                    5�_�   �   �           �   U   :    ����                                                                                                                                                                                                                                                                                                                            U          U          v       e���     �   T   V   �      R    getSum1Complement: somador port map (A => chOut, B => kpw, S => chComplement);5��    T   :                 �                    �    T   >                  �                     �    T   =                  �                     �    T   <                  �                     �    T   ;                  �                     �    T   :                 �                    �    T   :                 �                    �    T   :                 �                    5�_�   �   �           �   U   M    ����                                                                                                                                                                                                                                                                                                                            U          U          v       e���     �   T   V   �      [    getSum1Complement: somador port map (A => chOut, B => chComplement, S => chComplement);5��    T   M                 �                    �    T   R                  �                     �    T   Q                  �                     �    T   P                  �                     �    T   O                  �                     �    T   N                  �                     �    T   M                 �                    �    T   M                 �                    �    T   M                 �                    5�_�   �   �           �   U   Z    ����                                                                                                                                                                                                                                                                                                                            U          U          v       e���     �   U   W   �    �   U   V   �    5��    U                      �              ^       5�_�   �   �           �   V       ����                                                                                                                                                                                                                                                                                                                            V          V   
       v   
    e���     �   U   W   �      ]    getSum1Complement: somador port map (A => chOut, B => chComplement, S => sum1Complement);5��    U                     �                     5�_�   �   �           �   S   *    ����                                                                                                                                                                                                                                                                                                                            V          V   
       v   
    e��O     �   R   T   �      A    getE: somador port map (A => ei, B => sum1Out, S => preEOut);5��    R   *                 �
                    �    R   .                  �
                     �    R   -                  �
                     �    R   ,                  �
                     �    R   +                  �
                     �    R   *                 �
                    �    R   *                 �
                    �    R   *                 �
                    5�_�   �   �           �   S   F    ����                                                                                                                                                                                                                                                                                                                            V          V   
       v   
    e��f     �   R   S          G    getE: somador port map (A => ei, B => majComplement, S => preEOut);5��    R                      �
      H               5�_�   �   �           �   U   I    ����                                                                                                                                                                                                                                                                                                                            U          U   
       v   
    e��i     �   U   W   �    �   U   V   �    5��    U                      �              H       5�_�   �   �           �   U       ����                                                                                                                                                                                                                                                                                                                            U          U   
       v   
    e��q     �   T   V   �      Y    getComplement: somador port map (A => chOut, B => chComplement, S => sum1Complement);5��    T                     j                     5�_�   �   �           �   U   -    ����                                                                                                                                                                                                                                                                                                                            U          U   
       v   
    e���     �   T   V   �      \    getMajComplement: somador port map (A => chOut, B => chComplement, S => sum1Complement);5��    T   -                 �                    �    T   1                  �                     �    T   0                  �                     �    T   /                  �                     �    T   .                  �                     �    T   -                 �                    �    T   -                 �                    �    T   -                 �                    5�_�   �   �           �   U   N    ����                                                                                                                                                                                                                                                                                                                            U   N       U   Q       v   Q    e���     �   T   V   �      ^    getMajComplement: somador port map (A => sum1Out, B => chComplement, S => sum1Complement);5��    T   N                 �                    5�_�   �   �           �   V   F    ����                                                                                                                                                                                                                                                                                                                            U   N       U   Q       v   Q    e���     �   V   X   �    �   V   W   �    5��    V                      	              ^       5�_�   �   �   �       �   W       ����                                                                                                                                                                                                                                                                                                                            W          W   	       v   	    e���     �   V   X   �      ]    getMajComplement: somador port map (A => sum1Out, B => chComplement, S => majComplement);5��    V                                        5�_�   �   �           �   W   1    ����                                                                                                                                                                                                                                                                                                                            W          W   	       v   	    e���     �   V   X   �      ^    getSum0Complement: somador port map (A => sum1Out, B => chComplement, S => majComplement);5��    V   1                 :                    5�_�   �   �           �   W   <    ����                                                                                                                                                                                                                                                                                                                            W          W   	       v   	    e���     �   V   X   �      ^    getSum0Complement: somador port map (A => sum0Out, B => chComplement, S => majComplement);5��    V   <                 E                    �    V   A                  J                     �    V   @                  I                     �    V   ?                  H                     �    V   >                  G                     �    V   =                  F                     �    V   <                 E                    �    V   <                 E                    �    V   <                 E                    5�_�   �   �           �   W   Q    ����                                                                                                                                                                                                                                                                                                                            W          W   	       v   	    e���     �   V   X   �      `    getSum0Complement: somador port map (A => sum0Out, B => sum0Complement, S => majComplement);5��    V   Q                 Z                    �    V   T                  ]                     �    V   S                  \                     �    V   R                  [                     �    V   Q                 Z                    �    V   Q                 Z                    �    V   Q                 Z                    5�_�   �   �           �   Y        ����                                                                                                                                                                                                                                                                                                                            Y          h           V   W    e���     �   X   Y              -- Somadores       M    convertedIn1 <= signed('0' & di); -- extensão de sinal: número positivo   M    convertedIn2 <= signed('0' & hi); -- extensão de sinal: número positivo   N    convertedIn3 <= signed('0' & kpw); -- extensão de sinal: número positivo   R    convertedIn4 <= signed('0' & sum1_01); -- extensão de sinal: número positivo   O    convertedIn5 <= signed('0' & cho1); -- extensão de sinal: número positivo   R    convertedIn6 <= signed('0' & sum0_01); -- extensão de sinal: número positivo   O    convertedIn7 <= signed('0' & maj1); -- extensão de sinal: número positivo       Z    internal1 <= convertedIn1 + convertedIn2 + convertedIn3 + convertedIn4 + convertedIn5;   i    internal2 <= convertedIn2 + convertedIn3 + convertedIn4 + convertedIn5 + convertedIn6 + convertedIn7;       %    preOut1 <= bit_vector(internal1);   %    preOut2 <= bit_vector(internal2);    5��    X                      e      W              5�_�   �   �           �   Y       ����                                                                                                                                                                                                                                                                                                                            Y          Y           V   W    e���     �   X   Z   v          ao <= preOut2(31 downto 0);5��    X                     v                     5�_�   �   �           �   Y   
    ����                                                                                                                                                                                                                                                                                                                            Y          Y           V   W    e���     �   X   Z   v          ao <= preOut2;5��    X   
                 o                    �    X                    q                    �    X                     r                     �    X                     q                     �    X                     p                     �    X   
                 o                    �    X   
                 o                    �    X   
                 o                    5�_�   �   �           �   a       ����                                                                                                                                                                                                                                                                                                                            Y          Y           V   W    e���     �   `   b   v      
end arch7;5��    `                    �                    �    `                     �                     �    `                     �                     �    `                     �                     �    `                 
   �             
       �    `          
          �      
              �    `                 
   �             
       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            Y          Y           V   W    e���     �         v       architecture arch7 of stepfun is5��                                            �                     
                
       �              
                
              �                     
                
       5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                 V       e���     �             	   P    signal convertedIn1: signed(32 downto 0); -- entrada convertida para 33 bits   P    signal convertedIn2: signed(32 downto 0); -- entrada convertida para 33 bits   P    signal convertedIn3: signed(32 downto 0); -- entrada convertida para 33 bits   P    signal convertedIn4: signed(32 downto 0); -- entrada convertida para 33 bits   P    signal convertedIn5: signed(32 downto 0); -- entrada convertida para 33 bits   P    signal convertedIn6: signed(32 downto 0); -- entrada convertida para 33 bits   P    signal convertedIn7: signed(32 downto 0); -- entrada convertida para 33 bits   P    signal convertedIn8: signed(32 downto 0); -- entrada convertida para 33 bits    5��           	               3      �              5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                 V       e���     �                J    signal internal1: signed(32 downto 0);     -- somador interno: 33 bits   J    signal internal2: signed(32 downto 0);     -- somador interno: 33 bits5��                          �      �               5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                 V       e���     �         l          �         k    5��                          �                     �                         �                     5�_�   �   �           �      ,    ����                                                                                                                                                                                                                                                                                                                                                 V       e���     �         l      >    signal preAOut: bit_vector(31 downto 0);  -- pré-saida ao5��       ,                  :                     5�_�   �   �           �      ,    ����                                                                                                                                                                                                                                                                                                                                                 V       e���     �         l      >    signal preEOut: bit_vector(31 downto 0);  -- pré-saida eo5��       ,                  g                     5�_�   �   �           �   F       ����                                                                                                                                                                                                                                                                                                                                                 V       e��"     �   E   G   l      '    third: sum1 port map (ei, sum0Out);5��    E                    Q                    5�_�   �   �           �   G       ����                                                                                                                                                                                                                                                                                                                                                 V       e��#     �   F   H   l      (    fourth: sum0 port map (ai, sum1Out);5��    F                    z                    5�_�   �   �           �   G       ����                                                                                                                                                                                                                                                                                                                                                 V       e��0     �   F   H   l      (    fourth: sum1 port map (ai, sum1Out);5��    F                    �                    5�_�   �   �           �   F       ����                                                                                                                                                                                                                                                                                                                                                 V       e��6     �   E   G   l      '    third: sum0 port map (ei, sum0Out);5��    E                    ]                    5�_�   �   �           �   F       ����                                                                                                                                                                                                                                                                                                                                                 V       e��9    �   E   G   l      '    third: sum0 port map (1i, sum0Out);5��    E                    ]                    5�_�   �   �           �   L   !    ����                                                                                                                                                                                                                                                                                                                                                 V       e��y    �   K   M   l      G    getE: somador port map (A => ei, B => majComplement, S => preEOut);5��    K   !                 �                    5�_�   �   �           �   g        ����                                                                                                                                                                                                                                                                                                                                                 V       e���     �   f   g          T        carry(i+1) <= (A(i) and B(i)) or (A(i) and carry(i)) or (B(i) and carry(i));5��    f                      ;      U               5�_�   �   �           �   f        ����                                                                                                                                                                                                                                                                                                                                                 V       e���   	 �   e   g   k    �   f   g   k    5��    e                                    U       5�_�   �   �   �       �   f       ����                                                                                                                                                                                                                                                                                                                                                 V       e��Z     �   e   f          T        carry(i+1) <= (A(i) and B(i)) or (A(i) and carry(i)) or (B(i) and carry(i));5��    e                            U               5�_�   �   �           �   f       ����                                                                                                                                                                                                                                                                                                                                                 V       e��Z     �   f   h   k    �   f   g   k    5��    f                      ;              U       5�_�   �   �           �   D       ����                                                                                                                                                                                                                                                                                                                                                 V       e���     �   C   E   l      +    first: ch port map (ei, fi, gi, chOut);5��    C                    �                    5�_�   �   �           �   E       ����                                                                                                                                                                                                                                                                                                                                                 V       e���     �   D   F   l      .    second: maj port map (ai, bi, ci, majOut);5��    D                                        5�_�   �   �           �   E   	    ����                                                                                                                                                                                                                                                                                                                                                 V       e���     �   D   F   l      .    getMak: maj port map (ai, bi, ci, majOut);5��    D   	                                     5�_�   �   �           �   F       ����                                                                                                                                                                                                                                                                                                                                                 V       e���     �   E   G   l      '    third: sum0 port map (ai, sum0Out);5��    E                    G                    �    E                     N                     �    E   
                 M                    5�_�   �   �           �   G       ����                                                                                                                                                                                                                                                                                                                                                 V       e���    �   F   H   l      (    fourth: sum1 port map (ei, sum1Out);5��    F                    q                    5�_�   �   �   �       �           ����                                                                                                                                                                                                                                                                                                                               	       l   	       V   	    e��!     �         l       �         l    5��                         (               6       5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                               	       m   	       V   	    e��#     �         m    5��                          _                      5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                               	       n   	       V   	    e��%    �                use ieee.numeric_bit.all;5��                                                5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                               	       m   	       V   	    e��C     �         m      -- Declaração dos componentes5��                          �                     5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       e��E     �                 #    -- Declaração dos componentes�         n      #    -- Declaração dos componentes�      !   m    5��                        �      $       �      �                         �                    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       e��F     �                '        -- Declaração dos componentes�          n      '        -- Declaração dos componentes�         m    5��                        �      (       �      �                         �                    5�_�   �              �           ����                                                                                                                                                                                                                                                                                                                                      B           V       e��J     �             %   #    -- Declaração dos componentes       component ch is           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component maj is           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component sum0 is           port (   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component sum1 is           port (   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component somador is           port (   +            A : in bit_vector(31 downto 0);   +            B : in bit_vector(31 downto 0);   +            S : out bit_vector(31 downto 0)   
        );       end component;    5��           %               �      `              5�_�   �                       ����                                                                                                                                                                                                                                                                                                                                                 V       e��N     �         H    5��                          P                     �                          P                     �                          P                     5�_�                          ����                                                                                                                                                                                                                                                                                                                                                 V       e��O     �      3   I    �         I    5��                   %       P              `      5�_�                 3        ����                                                                                                                                                                                                                                                                                                                            D          D           V       e��S     �   2   3           5��    2                      �                     5�_�                 1       ����                                                                                                                                                                                                                                                                                                                            C          C           V       e��W     �   1   4   n          �   1   3   m    5��    1                      �                     �    1                      �                     �    1                     �                     �    2                  	   �              	       5�_�                 N   ;    ����                                                                                                                                                                                                                                                                                                                            E          E           V       e��z     �   M   O   o      ]    getMajComplement: somador port map (A => sum1Out, B => chComplement, S => majComplement);5��    M   ;                 �                    �    M   ?                  �                     �    M   >                  �                     �    M   =                  �                     �    M   <                  �                     �    M   ;                 �                    �    M   ;                 �                    �    M   ;                 �                    5�_�               P   <    ����                                                                                                                                                                                                                                                                                                                            E          E           V       e�Ǫ     �   P   R   o    �   P   Q   o    5��    P                      w	              H       5�_�                 Q       ����                                                                                                                                                                                                                                                                                                                            E          E           V       e�Ǭ     �   P   R   p      G    getE: somador port map (A => di, B => majComplement, S => preEOut);5��    P                    ~	                    5�_�    	             P   .    ����                                                                                                                                                                                                                                                                                                                            E          E           V       e�Ǹ     �   O   Q   p      Z    getSum0Complement: somador port map (A => sum0Out, B => sum0Complement, S => preAOut);5��    O   .                 J	                    �    O   1                  M	                     �    O   0                  L	                     �    O   /                  K	                     �    O   .                 J	                    �    O   .                 J	                    �    O   .                 J	                    5�_�    
          	   P   ;    ����                                                                                                                                                                                                                                                                                                                            E          E           V       e�Ǽ     �   O   Q   p      Y    getSum0Complement: somador port map (A => majOut, B => sum0Complement, S => preAOut);5��    O   ;                 W	                    �    O   @                  \	                     �    O   ?                  [	                     �    O   >                  Z	                     �    O   =                  Y	                     �    O   <                  X	                     �    O   ;                 W	                    �    O   ;                 W	                    �    O   ;                 W	                    5�_�  	            
   P   O    ����                                                                                                                                                                                                                                                                                                                            E          E           V       e���     �   O   Q   p      X    getSum0Complement: somador port map (A => majOut, B => majComplement, S => preAOut);5��    O   O                 k	                    �    O   T                  p	                     �    O   S                  o	                     �    O   R                  n	                     �    O   Q                  m	                     �    O   P                  l	                     �    O   O                 k	                    �    O   O                 k	                    �    O   O                 k	                    5�_�  
               Q   !    ����                                                                                                                                                                                                                                                                                                                            E          E           V       e���     �   P   R   p      G    getA: somador port map (A => di, B => majComplement, S => preEOut);5��    P   !                 �	                    �    P   %                  �	                     �    P   $                  �	                     �    P   #                  �	                     �    P   "                  �	                     �    P   !                 �	                    �    P   !                 �	                    �    P   !                 �	                    5�_�                 Q   /    ����                                                                                                                                                                                                                                                                                                                            E          E           V       e���     �   P   R   p      L    getA: somador port map (A => sum0Out, B => majComplement, S => preEOut);5��    P   /                 �	                    �    P   4                  �	                     �    P   3                  �	                     �    P   2                  �	                     �    P   1                  �	                     �    P   0                  �	                     �    P   /                 �	                    �    P   /                 �	                    �    P   /                 �	                    5�_�                 Q   G    ����                                                                                                                                                                                                                                                                                                                            E          E           V       e���    �   P   R   p      M    getA: somador port map (A => sum0Out, B => sum0Complement, S => preEOut);5��    P   G                 �	                    5�_�                   h       ����                                                                                                                                                                                                                                                                                                                            E          E           V       e���    �   g   h              carry(0) <= '0';5��    g                      _                     5�_�                 P   <    ����                                                                                                                                                                                                                                                                                                                            E          E           V       e�ǥ     �   P   Q   o    �   P   Q   o      Z    getSum0Complement: somador port map (A => sum0Out, B => sum0Complement, S => preAOut);5��    P                      w	              [       5�_�   �       �   �   �          ����                                                                                                                                                                                                                                                                                                                               	       m   	       V   	    e��     �         l    �         l      )use ieee.numeuse IEEE.STD_LOGIC_1164.ALL;   %use IEEE.NUMERIC_STD.ALL;ric_bit.all;5��                                       6       5�_�   �   �       �   �   D   
    ����                                                                                                                                                                                                                                                                                                                                                 V       e���     �   C   E        5��    C                      �      ,               5�_�   �   �           �   H   
    ����                                                                                                                                                                                                                                                                                                                                                 V       e���     �   H   I   k    �   H   I   k      +    getCh: ch port map (ei, fi, gi, chOut);5��    H                      �              ,       5�_�   �   �           �   F        ����                                                                                                                                                                                                                                                                                                                                                 V       e���     �   E   G        5��    E                      A      *               5�_�   �   �           �   I        ����                                                                                                                                                                                                                                                                                                                                                 V       e���     �   I   J   k    �   I   J   k      )    getSum1: sum1 port map (ei, sum1Out);5��    I                                    *       5�_�   �   �           �   D       ����                                                                                                                                                                                                                                                                                                                                                 V       e��3     �   C   E        5��    C                      �      /               5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                                                 V       e��4     �   K   L   k    �   K   L   k      .    getMaj: maj port map (ai, bi, ci, majOut);5��    K                      �              /       5�_�   �   �           �   D       ����                                                                                                                                                                                                                                                                                                                                                 V       e��:     �   C   E        5��    C                      �      *               5�_�   �   �           �   K        ����                                                                                                                                                                                                                                                                                                                                                 V       e��<    �   K   L   k    �   K   L   k      )    getSum0: sum0 port map (ai, sum0Out);5��    K                      �              *       5�_�   �               �   D        ����                                                                                                                                                                                                                                                                                                                                                 V       e��[    �   C   E        5��    C                      �                     5�_�   �           �   �   d       ����                                                                                                                                                                                                                                                                                                                                                 V       e��   
 �   c   e        5��    c                      �
                     5�_�   �           �   �   W       ����                                                                                                                                                                                                                                                                                                                            U   N       U   Q       v   Q    e���     �   V   X   �      ]    getlajComplement: somador port map (A => sum1Out, B => chComplement, S => majComplement);5��    V                                        5�_�   �           �   �   J       ����                                                                                                                                                                                                                                                                                                                            J          J   	       v       e��     �   J   K   {    �   J   K   {      '    third: sum1 port map (ei, sum1_01);5��    J                      �	              (       5�_�   y           {   z          ����                                                                                                                                                                                                                                                                                                                            ;          =                 e���     �         w    �         w      O    signal majOutchOut: signed(32 downto 0); -- entrada convertida para 33 bits5��                                              5�_�   P       Q   S   R   g       ����                                                                                                                                                                                                                                                                                                                            d          d          v       e�!     �   f   h   p      0    carry(0) <= '';  -- inicialização do carry5��    f                     �                     5�_�   P           R   Q   g       ����                                                                                                                                                                                                                                                                                                                            d          d          v       e� �     �   f   h        5��    f                      �      2               5�_�   @           B   A   _   &    ����                                                                                                                                                                                                                                                                                                                            \   
       \          v       e�g     �   ^   `   a      %        A: in bit_vector(31 downto 0)5��    ^   %                  �                     5�_�   6           8   7           ����                                                                                                                                                                                                                                                                                                                                                  V        e�     �       !   S    �       !   S          component maj is           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;    5��                           �              �       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �       F        5��            E                       �              5�_�                   M        ����                                                                                                                                                                                                                                                                                                                            C           E           V        e���     �   M   N   �    �   M   N   �      library ieee;   use ieee.numeric_bit.all;    5��    M                      �              )       5�_�                    M        ����                                                                                                                                                                                                                                                                                                                                                  V        e���     �   M   N   �    �   L   N   �      )5��    L                      �                     5�_�                    M        ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �   M   N   �    �   M   N   �      library ieee;   use ieee.numeric_bit.all;    5��    M                      �              )       5�_�                    .        ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �   .   /   �    �   .   /   �      library ieee;   use ieee.numeric_bit.all;    5��    .                      =              )       5�_�   	              
   #        ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �   #   $   �    �   #   $   �      library ieee;   use ieee.numeric_bit.all;    5��    #                      �              )       5�_�                    F       ����                                                                                                                                                                                                                                                                                                                                                             e���     �   E   G   �      O    signal convertedIn1: sined(32 downto 0); -- entrada convertida para 33 bits5��    E                     p                     5�_�                     F       ����                                                                                                                                                                                                                                                                                                                                                             e���     �   F   G   �    �   E   G   �      P    signal convertedIn1: singed(32 downto 0); -- entrada convertida para 33 bits5��    E                     q                     5��