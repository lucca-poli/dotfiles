Vim�UnDo� jo����f��
�\wksnH!�C���L�`   �                                  f=0    _�                             ����                                                                                                                                                                                                                                                                                                                                                             f=	}     �          �    �         �    5��                                           )       5�_�                    U       ����                                                                                                                                                                                                                                                                                                                                                             f=	�     �   T   V   �              if (clk'event) then5��    T          	          %      	              5�_�                    U       ����                                                                                                                                                                                                                                                                                                                                                             f=	�    �   T   V   �              if (clk) then5��    T                     $                     5�_�                    M       ����                                                                                                                                                                                                                                                                                                                                                             f=    �               �   library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity multisteps is   
    port (           clk, rst : in bit;   +        msgi : in bit_vector(511 downto 0);   -        haso : out bit_vector (255 downto 0);           done : out bit       );   end entity;       -architecture arch_multisteps of multisteps is       component stepfun is           port (   U                ai , bi , ci , di , ei , fi , gi , hi : in bit_vector (31 downto 0 );   2                kpw : in bit_vector (31 downto 0);   T                ao , bo , co , do , eo , fo , go , ho : out bit_vector (31 downto 0)   
        );       end component;              component somador is            port (   .            x, y: in bit_vector(31 downto 0);    *            q: out bit_vector(31 downto 0)           );        end component;           component sigma0 is            port(   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component sigma1 is           port(   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;       A    type wordArray is array (0 to 63) of bit_vector(31 downto 0);   @    type hashArray is array (0 to 7) of bit_vector(31 downto 0);       �    signal H : hashArray  := (X"6a09e667", X"bb67ae85", X"3c6ef372", X"a54ff53a", X"510e527f", X"9b05688c", X"1f83d9ab", X"5be0cd19");   �    signal K : wordArray := (X"428a2f98", X"71374491", X"b5c0fbcf", X"e9b5dba5", X"3956c25b", X"59f111f1", X"923f82a4", X"ab1c5ed5",   �                            X"d807aa98", X"12835b01", X"243185be", X"550c7dc3", X"72be5d74", X"80deb1fe", X"9bdc06a7", X"c19bf174",   �                            X"e49b69c1", X"efbe4786", X"0fc19dc6", X"240ca1cc", X"2de92c6f", X"4a7484aa", X"5cb0a9dc", X"76f988da",   �                            X"983e5152", X"a831c66d", X"b00327c8", X"bf597fc7", X"c6e00bf3", X"d5a79147", X"06ca6351", X"14292967",   �                            X"27b70a85", X"2e1b2138", X"4d2c6dfc", X"53380d13", X"650a7354", X"766a0abb", X"81c2c92e", X"92722c85",   �                            X"a2bfe8a1", X"a81a664b", X"c24b8b70", X"c76c51a3", X"d192e819", X"d6990624", X"f40e3585", X"106aa070",   �                            X"19a4c116", X"1e376c08", X"2748774c", X"34b0bcb5", X"391c0cb3", X"4ed8aa4a", X"5b9cca4f", X"682e6ff3",   �                            X"748f82ee", X"78a5636f", X"84c87814", X"8cc70208", X"90befffa", X"a4506ceb", X"bef9a3f7", X"c67178f2");       signal W, kpw : wordArray;   �    signal ain, bin, cin, din, ein, fin, gin, hin, kpwin, aout, bout, cout, dout, eout, fout, gout, hout: bit_vector(31 downto 0);       begin   $    w1_15: for i in 0 to 15 generate   	    begin   0        W(i) <= msgi((32*i + 31) downto (32*i));       end generate;       &    w16_63: for i in 16 to 63 generate   7    signal s1, s2, s3, s4, s5: bit_vector(31 downto 0);   	    begin   +        Soma1: sigma1 port map(W(i-2), s1);   ,        Soma2: sigma0 port map(W(i-15), s2);   0        Soma3: somador port map(s1, W(i-7), s3);   ,        Soma4: somador port map(s3, s2, s4);   1        Soma5: somador port map(s4, W(i-16), s5);           W(i) <= s5;       end generate;          (    kpw0_63: for j in 0 to 63 generate     	    begin   6        kpwsoma: somador port map(W(j), K(j), kpw(j));       end generate;          {    STEP: stepfun port map (ain, bin, cin, din, ein, fin, gin, hin, kpwin, aout, bout, cout, dout, eout, fout, gout, hout);           process(clk)       variable iterator: integer;   	    begin            if rising_edge(clk) then               if (rst = '1') then                   iterator := 0;                   done <= '0';       %            elsif (iterator = 0) then                   ain <= H(0);                   bin <= H(1);                   cin <= H(2);                   din <= H(3);   #                ein <= H(4);                          fin <= H(5);                   gin <= H(6);                   hin <= H(7);                    kpwin <= KPW(0);   )                iterator := iterator + 1;       &            elsif (iterator < 64) then                   ain <= aout;                   bin <= bout;                   cin <= cout;                   din <= dout;                   ein <= eout;                   fin <= fout;                   gin <= gout;                   hin <= hout;   '                kpwin <= KPW(iterator);   )                iterator := iterator + 1;                   else                   done <= '1';               end if;           end if;   end process;        =    SOMAF1: somador port map (aout, H(0), haso(31 downto 0));   >    SOMAF2: somador port map (bout, H(1), haso(63 downto 32));   >    SOMAF3: somador port map (cout, H(2), haso(95 downto 64));   ?    SOMAF4: somador port map (dout, H(3), haso(127 downto 96));   @    SOMAF5: somador port map (eout, H(4), haso(159 downto 128));   @    SOMAF6: somador port map (fout, H(5), haso(191 downto 160));   @    SOMAF7: somador port map (gout, H(6), haso(223 downto 192));   @    SOMAF8: somador port map (hout, H(7), haso(255 downto 224));       end architecture;       entity soma is   
    port (           a, b, carry: in bit;           sum, cout: out bit       );   end entity soma;        architecture ArchSoma of soma is   begin       sum <= (a xor b xor carry);   8    cout <= (a and b) or (a and carry) or (b and carry);        end architecture ArchSoma;       entity somador is   
    port (   *        x, y: in  bit_vector(31 downto 0);   '        q: out  bit_vector(31 downto 0)       );   end entity somador;       $architecture Archadder of somador is       component soma is           port (                a, b, carry: in bit;               sum, cout: out bit   
        );       end component;       (    signal aux: bit_vector(31 downto 0);   begin   9    SOMA0:  soma port map(x(0), y(0), '0', q(0), aux(0));   <    SOMA1:  soma port map(x(1), y(1), aux(0), q(1), aux(1));   <    SOMA2:  soma port map(x(2), y(2), aux(1), q(2), aux(2));   <    SOMA3:  soma port map(x(3), y(3), aux(2), q(3), aux(3));   <    SOMA4:  soma port map(x(4), y(4), aux(3), q(4), aux(4));   <    SOMA5:  soma port map(x(5), y(5), aux(4), q(5), aux(5));   <    SOMA6:  soma port map(x(6), y(6), aux(5), q(6), aux(6));   <    SOMA7:  soma port map(x(7), y(7), aux(6), q(7), aux(7));   <    SOMA8:  soma port map(x(8), y(8), aux(7), q(8), aux(8));   <    SOMA9:  soma port map(x(9), y(9), aux(8), q(9), aux(9));   @    SOMA10: soma port map(x(10), y(10), aux(9), q(10), aux(10));   A    SOMA11: soma port map(x(11), y(11), aux(10), q(11), aux(11));   A    SOMA12: soma port map(x(12), y(12), aux(11), q(12), aux(12));   A    SOMA13: soma port map(x(13), y(13), aux(12), q(13), aux(13));   A    SOMA14: soma port map(x(14), y(14), aux(13), q(14), aux(14));   A    SOMA15: soma port map(x(15), y(15), aux(14), q(15), aux(15));   A    SOMA16: soma port map(x(16), y(16), aux(15), q(16), aux(16));   A    SOMA17: soma port map(x(17), y(17), aux(16), q(17), aux(17));   A    SOMA18: soma port map(x(18), y(18), aux(17), q(18), aux(18));   A    SOMA19: soma port map(x(19), y(19), aux(18), q(19), aux(19));   A    SOMA20: soma port map(x(20), y(20), aux(19), q(20), aux(20));   A    SOMA21: soma port map(x(21), y(21), aux(20), q(21), aux(21));   A    SOMA22: soma port map(x(22), y(22), aux(21), q(22), aux(22));   A    SOMA23: soma port map(x(23), y(23), aux(22), q(23), aux(23));   A    SOMA24: soma port map(x(24), y(24), aux(23), q(24), aux(24));   A    SOMA25: soma port map(x(25), y(25), aux(24), q(25), aux(25));   A    SOMA26: soma port map(x(26), y(26), aux(25), q(26), aux(26));   A    SOMA27: soma port map(x(27), y(27), aux(26), q(27), aux(27));   A    SOMA28: soma port map(x(28), y(28), aux(27), q(28), aux(28));   A    SOMA29: soma port map(x(29), y(29), aux(28), q(29), aux(29));   A    SOMA30: soma port map(x(30), y(30), aux(29), q(30), aux(30));   A    SOMA31: soma port map(x(31), y(31), aux(30), q(31), aux(31));       end architecture Archadder;5�5�_�                     I       ����                                                                                                                                                                                                                                                                                                                                                             f=/    �               �   library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity multisteps is   
    port (           clk, rst : in bit;   +        msgi : in bit_vector(511 downto 0);   -        haso : out bit_vector (255 downto 0);           done : out bit       );   end entity;       -architecture arch_multisteps of multisteps is       component stepfun is           port (   U                ai , bi , ci , di , ei , fi , gi , hi : in bit_vector (31 downto 0 );   2                kpw : in bit_vector (31 downto 0);   T                ao , bo , co , do , eo , fo , go , ho : out bit_vector (31 downto 0)   
        );       end component;              component somador is            port (   .            x, y: in bit_vector(31 downto 0);    *            q: out bit_vector(31 downto 0)           );        end component;           component sigma0 is            port(   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component sigma1 is           port(   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;       A    type wordArray is array (0 to 63) of bit_vector(31 downto 0);   @    type hashArray is array (0 to 7) of bit_vector(31 downto 0);       �    signal H : hashArray  := (X"6a09e667", X"bb67ae85", X"3c6ef372", X"a54ff53a", X"510e527f", X"9b05688c", X"1f83d9ab", X"5be0cd19");   �    signal K : wordArray := (X"428a2f98", X"71374491", X"b5c0fbcf", X"e9b5dba5", X"3956c25b", X"59f111f1", X"923f82a4", X"ab1c5ed5",   �                            X"d807aa98", X"12835b01", X"243185be", X"550c7dc3", X"72be5d74", X"80deb1fe", X"9bdc06a7", X"c19bf174",   �                            X"e49b69c1", X"efbe4786", X"0fc19dc6", X"240ca1cc", X"2de92c6f", X"4a7484aa", X"5cb0a9dc", X"76f988da",   �                            X"983e5152", X"a831c66d", X"b00327c8", X"bf597fc7", X"c6e00bf3", X"d5a79147", X"06ca6351", X"14292967",   �                            X"27b70a85", X"2e1b2138", X"4d2c6dfc", X"53380d13", X"650a7354", X"766a0abb", X"81c2c92e", X"92722c85",   �                            X"a2bfe8a1", X"a81a664b", X"c24b8b70", X"c76c51a3", X"d192e819", X"d6990624", X"f40e3585", X"106aa070",   �                            X"19a4c116", X"1e376c08", X"2748774c", X"34b0bcb5", X"391c0cb3", X"4ed8aa4a", X"5b9cca4f", X"682e6ff3",   �                            X"748f82ee", X"78a5636f", X"84c87814", X"8cc70208", X"90befffa", X"a4506ceb", X"bef9a3f7", X"c67178f2");       signal W, kpw : wordArray;   �    signal ain, bin, cin, din, ein, fin, gin, hin, kpwin, aout, bout, cout, dout, eout, fout, gout, hout: bit_vector(31 downto 0);       begin   $    w1_15: for i in 0 to 15 generate   	    begin   0        W(i) <= msgi((32*i + 31) downto (32*i));       end generate;       &    w16_63: for i in 16 to 63 generate   7    signal s1, s2, s3, s4, s5: bit_vector(31 downto 0);   	    begin   +        Soma1: sigma1 port map(W(i-2), s1);   ,        Soma2: sigma0 port map(W(i-15), s2);   0        Soma3: somador port map(s1, W(i-7), s3);   ,        Soma4: somador port map(s3, s2, s4);   1        Soma5: somador port map(s4, W(i-16), s5);           W(i) <= s5;       end generate;          (    kpw0_63: for j in 0 to 63 generate     	    begin   6        kpwsoma: somador port map(W(j), K(j), kpw(j));       end generate;          {    STEP: stepfun port map (ain, bin, cin, din, ein, fin, gin, hin, kpwin, aout, bout, cout, dout, eout, fout, gout, hout);           process(clk)       variable iterator: integer;   	    begin            if rising_edge(clk) then               if (rst = '1') then                   iterator := 0;                   done <= '0';       %            elsif (iterator = 0) then                   ain <= H(0);                   bin <= H(1);                   cin <= H(2);                   din <= H(3);   #                ein <= H(4);                          fin <= H(5);                   gin <= H(6);                   hin <= H(7);                    kpwin <= KPW(0);   )                iterator := iterator + 1;       &            elsif (iterator < 64) then                   ain <= aout;                   bin <= bout;                   cin <= cout;                   din <= dout;                   ein <= eout;                   fin <= fout;                   gin <= gout;                   hin <= hout;   '                kpwin <= KPW(iterator);   )                iterator := iterator + 1;                   else                   done <= '1';               end if;           end if;   end process;        =    SOMAF1: somador port map (aout, H(0), haso(31 downto 0));   >    SOMAF2: somador port map (bout, H(1), haso(63 downto 32));   >    SOMAF3: somador port map (cout, H(2), haso(95 downto 64));   ?    SOMAF4: somador port map (dout, H(3), haso(127 downto 96));   @    SOMAF5: somador port map (eout, H(4), haso(159 downto 128));   @    SOMAF6: somador port map (fout, H(5), haso(191 downto 160));   @    SOMAF7: somador port map (gout, H(6), haso(223 downto 192));   @    SOMAF8: somador port map (hout, H(7), haso(255 downto 224));       end architecture;       entity soma is   
    port (           a, b, carry: in bit;           sum, cout: out bit       );   end entity soma;        architecture ArchSoma of soma is   begin       sum <= (a xor b xor carry);   8    cout <= (a and b) or (a and carry) or (b and carry);        end architecture ArchSoma;       entity somador is   
    port (   *        x, y: in  bit_vector(31 downto 0);   '        q: out  bit_vector(31 downto 0)       );   end entity somador;       $architecture Archadder of somador is       component soma is           port (                a, b, carry: in bit;               sum, cout: out bit   
        );       end component;       (    signal aux: bit_vector(31 downto 0);   begin   9    SOMA0:  soma port map(x(0), y(0), '0', q(0), aux(0));   <    SOMA1:  soma port map(x(1), y(1), aux(0), q(1), aux(1));   <    SOMA2:  soma port map(x(2), y(2), aux(1), q(2), aux(2));   <    SOMA3:  soma port map(x(3), y(3), aux(2), q(3), aux(3));   <    SOMA4:  soma port map(x(4), y(4), aux(3), q(4), aux(4));   <    SOMA5:  soma port map(x(5), y(5), aux(4), q(5), aux(5));   <    SOMA6:  soma port map(x(6), y(6), aux(5), q(6), aux(6));   <    SOMA7:  soma port map(x(7), y(7), aux(6), q(7), aux(7));   <    SOMA8:  soma port map(x(8), y(8), aux(7), q(8), aux(8));   <    SOMA9:  soma port map(x(9), y(9), aux(8), q(9), aux(9));   @    SOMA10: soma port map(x(10), y(10), aux(9), q(10), aux(10));   A    SOMA11: soma port map(x(11), y(11), aux(10), q(11), aux(11));   A    SOMA12: soma port map(x(12), y(12), aux(11), q(12), aux(12));   A    SOMA13: soma port map(x(13), y(13), aux(12), q(13), aux(13));   A    SOMA14: soma port map(x(14), y(14), aux(13), q(14), aux(14));   A    SOMA15: soma port map(x(15), y(15), aux(14), q(15), aux(15));   A    SOMA16: soma port map(x(16), y(16), aux(15), q(16), aux(16));   A    SOMA17: soma port map(x(17), y(17), aux(16), q(17), aux(17));   A    SOMA18: soma port map(x(18), y(18), aux(17), q(18), aux(18));   A    SOMA19: soma port map(x(19), y(19), aux(18), q(19), aux(19));   A    SOMA20: soma port map(x(20), y(20), aux(19), q(20), aux(20));   A    SOMA21: soma port map(x(21), y(21), aux(20), q(21), aux(21));   A    SOMA22: soma port map(x(22), y(22), aux(21), q(22), aux(22));   A    SOMA23: soma port map(x(23), y(23), aux(22), q(23), aux(23));   A    SOMA24: soma port map(x(24), y(24), aux(23), q(24), aux(24));   A    SOMA25: soma port map(x(25), y(25), aux(24), q(25), aux(25));   A    SOMA26: soma port map(x(26), y(26), aux(25), q(26), aux(26));   A    SOMA27: soma port map(x(27), y(27), aux(26), q(27), aux(27));   A    SOMA28: soma port map(x(28), y(28), aux(27), q(28), aux(28));   A    SOMA29: soma port map(x(29), y(29), aux(28), q(29), aux(29));   A    SOMA30: soma port map(x(30), y(30), aux(29), q(30), aux(30));   A    SOMA31: soma port map(x(31), y(31), aux(30), q(31), aux(31));       end architecture Archadder;5�5��