Vim�UnDo� �~��
���;{���_��ެ�#�A/u0�cv
�   d   entity contador_cm is             	       	   	   	    fs-    _�                            ����                                                                                                                                                                                                                                                                                                                                                             fs6     �   T   V          		digito2 => digito2,�   S   U          		digito1 => digito1,�   R   T          		digito0 => digito0,�   L   N          $	contador_bcd: contador_bcd_3digitos�   4   6          %	end component contador_bcd_3digitos;�   1   3          -			digito2: out std_logic_vector(3 downto 0);�   0   2          -			digito1: out std_logic_vector(3 downto 0);�   /   1          -			digito0: out std_logic_vector(3 downto 0);�   )   +          #	component contador_bcd_3digitos is�                ,		digito2: out std_logic_vector(3 downto 0);�                ,		digito1: out std_logic_vector(3 downto 0);�         d      ,		digito0: out std_logic_vector(3 downto 0);5��                        �                     �                        �                     �                        #                    �    )                                        �    /                    q                    �    0                    �                    �    1                    �                    �    4                    '                    �    L                    �                    �    R                    �                    �    R   
                 �                    �    S                    �                    �    S   
                 �                    �    T                                        �    T   
                                     5�_�                    *       ����                                                                                                                                                                                                                                                                                                                                                             fsI     �   )   +   d       	component contador_bcd_3digs is5��    )                                          5�_�                    5        ����                                                                                                                                                                                                                                                                                                                                                             fsO    �   4   6   d      "	end component contador_bcd_3digs;5��    4                      )                     5�_�                    M   !    ����                                                                                                                                                                                                                                                                                                                                                             fsc     �   L   N   d      !	contador_bcd: contador_bcd_3digs5��    L                      �                     5�_�                    M   
    ����                                                                                                                                                                                                                                                                                                                                                             fsk    �   L   N   d       	contador_bcd: contador_bcd_3dig5��    L   
                 �                    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             fs�    �   <   >          	contador_de_clock: contador_m�   '   )          	end component contador_m;�         d      	component contador_m is5��              
          �      
              �    '          
          �      
              �    <          
          �      
              5�_�      	              *        ����                                                                                                                                                                                                                                                                                                                                                             fs�    �   L   N          !	contador_digs: contador_bcd_3dig�   4   6          !	end component contador_bcd_3dig;�   )   +   d      	component contador_bcd_3dig is5��    )                                        �    4                    "                    �    L                    �                    5�_�                  	           ����                                                                                                                                                                                                                                                                                                                                                             fs,    �   c   e          "end architecture contador_cm_arch;�                /architecture contador_cm_arch of contador_cm is�                end entity contador_cm;�         d      entity contador_cm is5��                        3                     �                        �                    �                        �                    �       $                 �                    �    c                    $                    5�_�                             ����                                                                                                                                                                                                                                                                                                                                                             fs-     �         d      )		gig0: out std_logic_vector(3 downto 0);�                )		gig1: out std_logic_vector(3 downto 0);�                )		gig2: out std_logic_vector(3 downto 0);�   )   +           	component contador_bcd_3gigs is�   /   1          *			gig0: out std_logic_vector(3 downto 0);�   0   2          *			gig1: out std_logic_vector(3 downto 0);�   1   3          *			gig2: out std_logic_vector(3 downto 0);�   4   6          "	end component contador_bcd_3gigs;�   L   N          !	contador_bcd: contador_bcd_3gigs�   R   T          		gig0 => digito0,�   S   U          		gig1 => digito1,�   T   V          		gig2 => digito2,5��                        �                     �                        �                     �                        #                    �    )                                        �    /                    q                    �    0                    �                    �    1                    �                    �    4                    '                    �    L                    �                    �    R                    �                    �    S                    �                    �    T                    
                    5��