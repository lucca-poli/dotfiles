Vim�UnDo� mc��aZȍ��)�p'��6�7!Q�]i���0   \   "use IEEE.NUMERIC_BIT_UNSIGNED.ALL;   #          _       _   _   _    e��    _�                           ����                                                                                                                                                                                                                                                                                                                                                             e�O     �         ^    �         ^    5��                                        G       5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �      
   b      +	signal op1, op2 : bit_vector(31 downto 0);5��                         �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �                    a <= x and y;5��                                               5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �         a          op2 <= ((not x) and z);5��                         �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �         a          op2 <= ((not x) and z;5��                         �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �                    b <= not(x) and z;5��                                               5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �                    c <= a xor b;5��                                               5�_�                       	    ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �         _          q <= c;5��       	                                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �         _          q <= op1 xor op2; 5��                        �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �         _      /	signal op1, op2, op3: bit_vector(31 downto 0);5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �      $   _    �         _    5��                          W              Z       5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �                     b <= x and z;5��                          i                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �                     c <= y and x;5��                          i                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �                    a <= z and y;5��                          W                     5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �         a          q <= op1 xor op2 xor op3; 5��                        <                    5�_�       "           !          ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �                    d <= a xor b xor c;5��                          Y                     5�_�   !   #           "      	    ����                                                                                                                                                                                                                                                                                                                                                             e�O�     �          `          q <= d;5��       	                 b                    5�_�   "   $           #   /       ����                                                                                                                                                                                                                                                                                                                                                             e�P�     �   /   1   `    �   /   0   `    5��    /                      V              2       5�_�   #   &           $   ,       ����                                                                                                                                                                                                                                                                                                                            /          ,          V       e�Q     �   +   ,          K	rot2 <= (31 downto 30 => x(1 downto 0)) & (29 downto 0 => x(31 downto 2));   Q    rot13 <= (31 downto 19 => x(12 downto 0)) & (18 downto 0 => x(31 downto 13));   P    rot22 <= (31 downto 10 => x(21 downto 0)) & (9 downto 0 => x(31 downto 22));   "    q <= rot2 xor rot13 xor rot22;5��    +                      D                    5�_�   $   '   %       &   *       ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       e�Q?     �   )   *          4	signal rot2, rot13, rot22: bit_vector(31 downto 0);5��    )                      	      5               5�_�   &   (           '   :       ����                                                                                                                                                                                                                                                                                                                            +          +          V       e�QO     �   :   <   \    �   :   ;   \    5��    :                                    6       5�_�   '   )           (   <       ����                                                                                                                                                                                                                                                                                                                            +          +          V       e�QQ     �   ;   <          "    q <= rot6 xor rot11 xor rot25;5��    ;                      B      #               5�_�   (   *           )   8       ����                                                                                                                                                                                                                                                                                                                            +          +          V       e�QZ     �   7   8          K	rot6 <= (31 downto 26 => x(5 downto 0)) & (25 downto 0 => x(31 downto 6));   Q    rot11 <= (31 downto 21 => x(10 downto 0)) & (20 downto 0 => x(31 downto 11));   O    rot25 <= (31 downto 7 => x(24 downto 0)) & (6 downto 0 => x(31 downto 25));5��    7                            �               5�_�   )   +           *   6       ����                                                                                                                                                                                                                                                                                                                            +          +          V       e�Q\     �   5   6          4	signal rot6, rot11, rot25: bit_vector(31 downto 0);5��    5                      �      5               5�_�   *   ,           +   7       ����                                                                                                                                                                                                                                                                                                                            +          +          V       e�Q]     �   6   8   X      5        q <= (x ror 6) xor (x ror 11) xor (x ror 25);5��    6                     �                     5�_�   +   -           ,   E        ����                                                                                                                                                                                                                                                                                                                            D           G          V       e�Qo     �   C   E   U      K	rot7 <= (31 downto 25 => x(6 downto 0)) & (24 downto 0 => x(31 downto 7));�   D   E          Q    rot18 <= (31 downto 14 => x(17 downto 0)) & (13 downto 0 => x(31 downto 18));   C    sr3 <= (31 downto 29 => '0') & (28 downto 0 => x(31 downto 3));        q <= rot7 xor rot18 xor sr3;5��    D                      H      �               �    C          J           �      J               �    C                     �                    �    C                      �                     5�_�   ,   .           -   D        ����                                                                                                                                                                                                                                                                                                                            D           E          V       e�Qp     �   D   I   U    �   D   E   U    5��    D                      �                    5�_�   -   /           .   D        ����                                                                                                                                                                                                                                                                                                                            D           I          V       e�Qq     �   C   D           5��    C                      �                     5�_�   .   0           /   D       ����                                                                                                                                                                                                                                                                                                                            D           H          V       e�Qu     �   C   D          K	rot7 <= (31 downto 25 => x(6 downto 0)) & (24 downto 0 => x(31 downto 7));   Q    rot18 <= (31 downto 14 => x(17 downto 0)) & (13 downto 0 => x(31 downto 18));   C    sr3 <= (31 downto 29 => '0') & (28 downto 0 => x(31 downto 3));        q <= rot7 xor rot18 xor sr3;5��    C                      �                    5�_�   /   1           0   D       ����                                                                                                                                                                                                                                                                                                                            D           D          V       e�Qy     �   C   E   T    �   D   E   T    5��    C                      �              5       5�_�   0   2           1   D       ����                                                                                                                                                                                                                                                                                                                            E           E          V       e�Qz     �   C   E   U      4        q <= (x ror 7) xor (x ror 18) xor (x srl 3);5��    C                                           5�_�   1   3           2   B        ����                                                                                                                                                                                                                                                                                                                            E           E          V       e�Q{     �   A   B          2	signal rot7, rot18, sr3: bit_vector(31 downto 0);5��    A                      �      3               5�_�   2   4           3   P        ����                                                                                                                                                                                                                                                                                                                            S          P           V       e�Q�     �   O   P          N	rot17 <= (31 downto 15 => x(16 downto 0)) & (14 downto 0 => x(31 downto 17));   Q    rot19 <= (31 downto 13 => x(18 downto 0)) & (12 downto 0 => x(31 downto 19));   E    sr10 <= (31 downto 22 => '0') & (21 downto 0 => x(31 downto 10));   "    q <= rot17 xor rot19 xor sr10;5��    O                      �      
              5�_�   3   5           4   N        ����                                                                                                                                                                                                                                                                                                                            P          P           V       e�Q�     �   M   N          4	signal rot17, rot19, sr10: bit_vector(31 downto 0);5��    M                      �      5               5�_�   4   6           5   N       ����                                                                                                                                                                                                                                                                                                                            O          O           V       e�Q�     �   N   P   O    �   N   O   O    5��    N                      �              7       5�_�   5   7           6   O       ����                                                                                                                                                                                                                                                                                                                            P          P           V       e�Q�    �   N   P   P      6        q <= (x ror 17) xor (x ror 19) xor (x srl 10);5��    N                     �                     5�_�   6   8           7          ����                                                                                                                                                                                                                                                                                                                                                V       e�Rj     �          P    �         P    5��                                           (       5�_�   7   9           8           ����                                                                                                                                                                                                                                                                                                                                                V       e�Rk   	 �         R    5��                          (                      5�_�   8   ;           9           ����                                                                                                                                                                                                                                                                                                                                       S           V        e�[x     �               S   library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity ch is   	port (   )    	x, y, z: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end ch;       architecture arch1 of ch is   0	signal op1, op2, op3 : bit_vector(31 downto 0);   begin   	op1 <= x and y;       op2 <= (not x) and z;       op3 <= op1 xor op2;        q <= op3;   
end arch1;       entity maj is   	port (   )    	x, y, z: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end maj;       architecture arch2 of maj is   4	signal op1, op2, op3, op4: bit_vector(31 downto 0);   begin   	op1 <= x and y;       op2 <= x and z;       op3 <= y and z;        op4 <= op1 xor op2 xor op3;        q <= op4;   
end arch2;       entity sum0 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   	end sum0;       architecture arch3 of sum0 is   begin   1    q <= (x ror 2) xor (x ror 13) xor (x ror 22);   
end arch3;       entity sum1 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   	end sum1;       architecture arch4 of sum1 is   begin   1    q <= (x ror 6) xor (x ror 11) xor (x ror 25);   
end arch4;       entity sigma0 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end sigma0;       architecture arch5 of sigma0 is   begin   0    q <= (x ror 7) xor (x ror 18) xor (x srl 3);   
end arch5;       entity sigma1 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end sigma1;       architecture arch6 of sigma1 is   begin   2    q <= (x ror 17) xor (x ror 19) xor (x srl 10);   
end arch6;5�5�_�   9   =   :       ;      	    ����                                                                                                                                                                                                                                                                                                                                                             e��     �         T      use IEEE.std_logic_1164.ALL;5��       	                 1                     �                         3                      �       
                 2                     �                         3                      �       
                  2                      �       	                 1                     �                         3                      �       
                  2                      �       	                 1                     �       	                 1                     �       	                 1                     �       	                 1                     �       	                 1                     5�_�   ;   ?   <       =   %        ����                                                                                                                                                                                                                                                                                                                                                  V        e��$     �   %   *   T    �   %   &   T    5��    %                      �              C       5�_�   =   @   >       ?   5        ����                                                                                                                                                                                                                                                                                                                                                  V        e��+     �   5   :   X    �   5   6   X    5��    5                      �              C       5�_�   ?   A           @   E        ����                                                                                                                                                                                                                                                                                                                                                  V        e��-     �   E   J   \    �   E   F   \    5��    E                      �              C       5�_�   @   C           A   U        ����                                                                                                                                                                                                                                                                                                                                                  V        e��0     �   U   Z   `    �   U   V   `    5��    U                                    C       5�_�   A   D   B       C   X   	    ����                                                                                                                                                                                                                                                                                                                                                  V        e��6     �   W   Y   d      use IEEE.NUMERIC_STD.ALL;5��    W   	                 C                    �    W                     E                     �    W   
                  D                     �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    5�_�   C   E           D   X   	    ����                                                                                                                                                                                                                                                                                                                                                  V        e��?     �   W   Y   d      "use IEEE.NUMERIC_BIT_UNSIGNED.ALL;5��    W   	                 C                    �    W                     F                     �    W                     E                     �    W   
                  D                     �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    5�_�   D   F           E   X   	    ����                                                                                                                                                                                                                                                                                                                                                  V        e��G     �   W   Y   d      "use IEEE.NUMERIC_STD_UNSIGNED.ALL;5��    W   	                 C                    �    W                     E                     �    W   
                  D                     �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    �    W   	                 C                    5�_�   E   G           F   H       ����                                                                                                                                                                                                                                                                                                                                                  V        e��S     �   H   J   d    �   H   I   d    5��    H                      2              #       5�_�   F   H           G   H        ����                                                                                                                                                                                                                                                                                                                                                  V        e��T     �   G   H          use IEEE.NUMERIC_STD.ALL;5��    G                                           5�_�   G   I           H   8        ����                                                                                                                                                                                                                                                                                                                                                  V        e��Z     �   8   :   d    �   8   9   d    5��    8                                    #       5�_�   H   J           I   8        ����                                                                                                                                                                                                                                                                                                                                                  V        e��[     �   7   8          use IEEE.NUMERIC_STD.ALL;5��    7                      �                     5�_�   I   K           J   (        ����                                                                                                                                                                                                                                                                                                                                                  V        e��^     �   (   *   d    �   (   )   d    5��    (                      �              #       5�_�   J   L           K   (        ����                                                                                                                                                                                                                                                                                                                                                  V        e��_   
 �   '   (          use IEEE.NUMERIC_STD.ALL;5��    '                      �                     5�_�   K   M           L   '        ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �   &   '          use IEEE.NUMERIC_BIT.ALL;5��    &                      �                     5�_�   L   N           M           ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �                use IEEE.NUMERIC_BIT.ALL;5��                                                5�_�   M   O           N   5        ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �   4   5          use IEEE.NUMERIC_BIT.ALL;5��    4                      �                     5�_�   N   P           O   D        ����                                                                                                                                                                                                                                                                                                                                                  V        e��     �   C   D          use IEEE.NUMERIC_BIT.ALL;5��    C                      �                     5�_�   O   Q           P   S        ����                                                                                                                                                                                                                                                                                                                                                  V        e��    �   R   S          use IEEE.NUMERIC_BIT.ALL;5��    R                      �                     5�_�   P   R           Q      	    ����                                                                                                                                                                                                                                                                                                                                                  V        e�     �                use IEEE.NUMERIC_STD.ALL;5��                                                5�_�   Q   S           R           ����                                                                                                                                                                                                                                                                                                                                                  V        e�     �                 library IEEE;5��                                                  5�_�   R   \           S           ����                                                                                                                                                                                                                                                                                                                                                  V        e�    �                  5��                                                  5�_�   S   ]   [       \   #   	    ����                                                                                                                                                                                                                                                                                                                            "   	       #   	       V   	    e��    �   !   $   \      library IEEE;   "use IEEE.NUMERIC_BIT_UNSIGNED.ALL;5��    !                     s      1       7       5�_�   \   ^           ]   2   	    ����                                                                                                                                                                                                                                                                                                                            1   	       2   	       V   	    e��     �   0   3   \      library IEEE;   "use IEEE.NUMERIC_BIT_UNSIGNED.ALL;5��    0                     �      1       7       5�_�   ]   _           ^   A   	    ����                                                                                                                                                                                                                                                                                                                            @   	       A   	       V   	    e��     �   ?   B   \      library IEEE;   "use IEEE.NUMERIC_BIT_UNSIGNED.ALL;5��    ?                     �      1       7       5�_�   ^               _   P   	    ����                                                                                                                                                                                                                                                                                                                            O   	       P   	       V   	    e��    �   N   Q   \      library IEEE;   "use IEEE.NUMERIC_BIT_UNSIGNED.ALL;5��    N                     �      1       7       5�_�   S       Y   \   [   O   	    ����                                                                                                                                                                                                                                                                                                                            P   	       O   	       V   	    e��     �   N   Q   \      -- library IEEE;   %-- use IEEE.NUMERIC_BIT_UNSIGNED.ALL;5��    N                     �      1       7       5�_�   S   Z   X   [   Y   A   	    ����                                                                                                                                                                                                                                                                                                                            /   	                 V       e�h    �   @   B   \      "use IEEE.NUMERIC_BIT_UNSIGNED.ALL;5��    @   	                 �                    �    @                     �                     �    @   
                  �                     �    @   	                 �                    �    @   	                 �                    �    @   	                 �                    �    @   	                 �                    �    @   	                 �                    �    @                     �                     �    @   
                  �                     �    @   	                 �                    �    @   	                 �                    �    @   	                 �                    �    @   	                 �                    5�_�   Y               Z   #        ����                                                                                                                                                                                                                                                                                                                            0   	                 V       e��     �   #   $   \    �   "   $   \      use IEEE.STD_LOGIC_1164.ALL;   use IEEE.NUMERIC_STD.ALL;5��    "           "           �      "               �    "                     �              6       5�_�   S       W   Y   X   O        ����                                                                                                                                                                                                                                                                                                                                                  V        e�(     �   N   R        5��    N                      �      2               5�_�   S       V   X   W   @        ����                                                                                                                                                                                                                                                                                                                                                  V        e�$     �   ?   C        5��    ?                      �      2               5�_�   S       U   W   V   1        ����                                                                                                                                                                                                                                                                                                                                                  V        e�      �   0   4        5��    0                            2               5�_�   S       T   V   U   1        ����                                                                                                                                                                                                                                                                                                                                                  V        e�     �   0   4        5��    0                            2               5�_�   S           U   T   "        ����                                                                                                                                                                                                                                                                                                                                                  V        e�     �   !   %        5��    !                      s      2               5�_�   A           C   B   X        ����                                                                                                                                                                                                                                                                                                                                                  V        e��4     �   W   Y        5��    W                      :                     5�_�   =           ?   >   0        ����                                                                                                                                                                                                                                                                                                                                                  V        e��(     �   0   1   X    �   0   1   X      library IEEE;   use IEEE.NUMERIC_BIT.ALL;   use IEEE.NUMERIC_STD.ALL;    5��    0                      q              C       5�_�   ;           =   <           ����                                                                                                                                                                                                                                                                                                                                                  V        e��!     �         T    �         T      library IEEE;   use IEEE.NUMERIC_BIT.ALL;   use IEEE.NUMERIC_STD.ALL;    5��                          �               C       5�_�   9           ;   :           ����                                                                                                                                                                                                                                                                                                                                                             e��     �              5��                          (                      5�_�   $           &   %   *       ����                                                                                                                                                                                                                                                                                                                            +          +          V       e�Q;     �   )   +        5��    )                      	      5               5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�O     �         ^          q <= op2 xor op2; 5��                                             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �      	   ^       architecture behavioral of ch is5��                     
   �              
       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �         ^      end behavioral;5��                                            �                                              �                                              �                     
                
       �              
                
              �                     
                
       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �         ^      architecture beh of maj is5��                        �                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �         ^      architecture beh[] of maj is5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �         ^      !architecture behavioral of maj is5��                         �                     �                     
   �             
       �              
          �      
              �                     
   �             
       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �         ^      end be;5��                        R                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �         ^      	end be[];5��                         T                     5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �         ^      end behavioral;5��                         T                     �                         T                     �                         S                     �                     
   R             
       �              
          R      
              �                     
   R             
       5�_�      
           	   '       ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �   &   (   ^      "architecture behavioral of sum0 is5��    &                    �                    �    &                 
   �             
       �    &          
          �      
              �    &                 
   �             
       5�_�   	              
   .       ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �   -   /   ^      end behavioral;5��    -                    K                    �    -                     L                     �    -                 
   K             
       �    -          
          K      
              �    -                 
   K             
       5�_�   
                 7       ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �   6   8   ^      "architecture behavioral of sum1 is5��    6                    �                    �    6                 
   �             
       �    6          
          �      
              �    6                 
   �             
       5�_�                    >       ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �   =   ?   ^      end behavioral;5��    =                    C                    �    =                     E                     �    =                     D                     �    =                 
   C             
       �    =          
          C      
              �    =                 
   C             
       5�_�                    G       ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �   F   H   ^      $architecture behavioral of sigma0 is5��    F                    �                    �    F                 
   �             
       �    F          
          �      
              �    F                 
   �             
       5�_�                    N       ����                                                                                                                                                                                                                                                                                                                                                             e�L      �   M   O   ^      end behavioral;5��    M                    1                    �    M                     2                     �    M                 
   1             
       �    M          
          1      
              �    M                 
   1             
       5�_�                    W       ����                                                                                                                                                                                                                                                                                                                                                             e�L     �   V   X   ^      $architecture behavioral of sigma1 is5��    V                    �                    �    V                 
   �             
       �    V          
          �      
              �    V                 
   �             
       5�_�                     ^       ����                                                                                                                                                                                                                                                                                                                                                             e�L    �   ]   _          end behavioral;5��    ]                    (
                    �    ]                     )
                     �    ]                 
   (
             
       �    ]          
          (
      
              �    ]                 
   (
             
       5��