Vim�UnDo� �B���;���$F�U�����d��j�h!   X   entity interface_hcsr04 is                              fs�    _�                              ����                                                                                                                                                                                                                                                                                                                                                             fs�    �   W   Y          'end architecture interface_hcsr04_arch;�   E   G          	UC: interface_hcsr04_uc�   7   9          	FD: interface_hcsr04_fd�   1   3          #	end component interface_hcsr04_uc;�   #   %          !	component interface_hcsr04_uc is�   !   #          #	end component interface_hcsr04_fd;�                !	component interface_hcsr04_fd is�                9architecture interface_hcsr04_arch of interface_hcsr04 is�                end entity interface_hcsr04;�         X      entity interface_hcsr04 is5��                        3                     �                        }                    �                        �                    �       %                 �                    �                        �                    �    !                    �                    �    #                                        �    1                    c                    �    7                    �                    �    E                    �                    �    W                    �                    5��