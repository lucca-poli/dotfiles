Vim�UnDo� 0ߠ��l��χ@\��Ԝ�a'z�%��@����   �   (    w_vec(0)  <= msgi(31 downto 0); -- 0   x   (                       f��    _�                             ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�'     �         '    5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�*     �         (    5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�+     �         )       �        )    5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�-     �                 antonio.seabra@usp.br5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�H     �         )       �        )    5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�I     �                 antonio.seabra@usp.br5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�P     �         )       �        )    5��                                           #      5�_�      	                      ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�Q     �                 5��                          #                     5�_�                 	           ����                                                                                                                                                                                                                                                                                                                                                 V       f�i    �                 library IEEE;   "use IEEE.NUMERIC_BIT_UNSIGNED.ALL;       entity sigma0 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end sigma0;       architecture arch5 of sigma0 is   begin   0    q <= (x ror 7) xor (x ror 18) xor (x srl 3);   
end arch5;       library IEEE;   "use IEEE.NUMERIC_BIT_UNSIGNED.ALL;       entity sigma1 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end sigma1;       architecture arch6 of sigma1 is   begin   2    q <= (x ror 17) xor (x ror 19) xor (x srl 10);   
end arch6;    5��                                   $              5�_�   	                        ����                                                                                                                                                                                                                                                                                                                            �   G       �   G       V   G    f6�    �  &  (          end somadorarch;�   �   �          &architecture somadorarch of somador is�   �   �          end somador;�   �   �          entity somador is�   �   �          	--somador�   �   �          ^        inst13: somador port map (a => hout, b => x"5be0cd19",  soma => haso(255 downto 224));�   �   �          ^        inst12: somador port map (a => gout, b => x"1f83d9ab",  soma => haso(223 downto 192));�   �   �          ^        inst11: somador port map (a => fout, b => x"9b05688c",  soma => haso(191 downto 160));�   �   �          ^        inst10: somador port map (a => eout, b => x"510e527f",  soma => haso(159 downto 128));�   �   �          \        inst9: somador port map (a => dout, b => x"a54ff53a",  soma => haso(127 downto 96));�   �   �          [        inst8: somador port map (a => cout, b => x"3c6ef372",  soma => haso(95 downto 64));�   �   �          [        inst7: somador port map (a => bout, b => x"bb67ae85",  soma => haso(63 downto 32));�   �   �          Z        inst6: somador port map (a => aout, b => x"6a09e667",  soma => haso(31 downto 0));�   �   �          E        	sum: somador port map(a => waux, b => kaux, soma => kpwaux);�   �   �          2        	inst5: somador port map(y4, W(i-16), y5);�   �   �          -        	inst4: somador port map(y3, y2, y4);�   �   �          1        	inst3: somador port map(y1, W(i-7), y3);�        '      component somador is5��       
              
   �             
       �    �                 
   �             
       �    �                 
   �             
       �    �                 
                
       �    �                 
                
       �    �                 
   �             
       �    �                 
                
       �    �                 
   x             
       �    �                 
   �             
       �    �                 
   8             
       �    �                 
   �             
       �    �                 
   �             
       �    �                 
   ^             
       �    �                 
   �             
       �    �                 
   �             
       �    �                 
   N             
       �    �                 
   h             
       �    �                 
   z             
       �    &                
   �'             
       5�_�                            ����                                                                                                                                                                                                                                                                                                                            �   G       �   G       V   G    f6�    �                +architecture arqmultisteps of multisteps is�        '      entity multisteps is5��              
          0       
              �              
          �       
              �       !       
                
              5�_�                    �   J    ����                                                                                                                                                                                                                                                                                                                            �   J       �   J          J    fYJ    �   �   �  '      ^        inst7: somador_v0 port map (a => bout, b => x"bb67ae85",  soma => haso(63 downto 32));   ^        inst8: somador_v0 port map (a => cout, b => x"3c6ef372",  soma => haso(95 downto 64));   _        inst9: somador_v0 port map (a => dout, b => x"a54ff53a",  soma => haso(127 downto 96));�   �   �  '      ]        inst6: somador_v0 port map (a => aout, b => x"6a09e667",  soma => haso(31 downto 0));5��    �   J                  �                     �    �   J                  ^                     �    �   J                  �                     �    �   J                                       5�_�                    2       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   1   2          Ksignal s1, s2, s3, s4, sa, sb, sc, sd, sW, se, sf: bit_vector(31 downto 0);5��    1                      �      L               5�_�                    4       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   3   4          signal step: integer; 5��    3                      �                     5�_�                    3   7    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   2   4  %      Wsignal aout, bout, cout, dout, eout, fout, gout, hout, kpwout: bit_vector(31 downto 0);5��    2   7                  `                     5�_�                    3   5    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   2   4  %      Qsignal aout, bout, cout, dout, eout, fout, gout, hout, : bit_vector(31 downto 0);5��    2   5                  ^                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �          &    soma : out bit_vector(31 downto 0)�   �   �          a        inst13: somador_v0 port map (a => hout, b => x"5be0cd19",  soma => haso(255 downto 224));�   �   �          a        inst12: somador_v0 port map (a => gout, b => x"1f83d9ab",  soma => haso(223 downto 192));�   �   �          a        inst11: somador_v0 port map (a => fout, b => x"9b05688c",  soma => haso(191 downto 160));�   �   �          a        inst10: somador_v0 port map (a => eout, b => x"510e527f",  soma => haso(159 downto 128));�   �   �          `        inst9: somador_v0 port map (a => dout, b => x"a54ff53a",  soma =>  haso(127 downto 96));�   �   �          _        inst8: somador_v0 port map (a => cout, b => x"3c6ef372",  soma =>  haso(95 downto 64));�   �   �          _        inst7: somador_v0 port map (a => bout, b => x"bb67ae85",  soma =>  haso(63 downto 32));�   �   �          ^        inst6: somador_v0 port map (a => aout, b => x"6a09e667",  soma =>  haso(31 downto 0));�   �   �          $                        hin <= hout;�   �   �          $                        gin <= gout;�   �   �          $                        fin <= fout;�   �   �          $                        ein <= eout;�   �   �          $                        din <= dout;�   �   �          $                        cin <= cout;�   �   �          $                        bin <= bout;�   �   �          $                        ain <= aout;�   �   �          t        inststep : stepfun port map (ain,bin,cin,din,ein,fin,gin,hin,kpwin,aout,bout,cout,dout,eout,fout,gout,hout);�   2   4          Osignal aout, bout, cout, dout, eout, fout, gout, hout: bit_vector(31 downto 0);�   (   *          &        q: out bit_vector(31 downto 0)�   !   #          &        q: out bit_vector(31 downto 0)�                &    soma : out bit_vector(31 downto 0)�                7  ao,bo,co,do,eo,fo,go,ho: out bit_vector (31 downto 0)�      
                  done : out bit�      	  %      ,        haso : out bit_vector(255 downto 0);5��                        �                     �                        �                     �                        �                    �                        7                    �    !                    �                    �    (                    A                    �    2                    7                    �    2                    >                    �    2                    E                    �    2                    L                    �    2   $                 S                    �    2   +                 Z                    �    2   2                 a                    �    2   9                 h                    �    �   L                 �                    �    �   R                 �                    �    �   X                 �                    �    �   ^                 �                    �    �   d                 �                    �    �   j                 �                    �    �   p                 �                    �    �   v                 �                    �    �                     �                    �    �                                         �    �                     <                    �    �                     b                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     �                    �    �   *                 �                    �    �   *                 �                    �    �   *                 S                    �    �   *                 �                    �    �   +                                     �    �   +                 z                    �    �   +                 �                    �    �   +                 @                    �    �                    �                    5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �  %      '    soma : _out bit_vector(31 downto 0)5��    �                     �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�      �      	  %      -        haso : _out bit_vector(255 downto 0);5��                         �                      5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                             f�     �      
  %              done : _out bit5��                         �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�     �        %      8  ao,bo,co,do,eo,fo,go,ho: _out bit_vector (31 downto 0)5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�     �        %      '    soma : _out bit_vector(31 downto 0)5��                         4                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�     �        %      &    soma : out bit_vector(31 downto 0)5��                        -                    5�_�                   %       ����                                                                                                                                                                                                                                                                                                                                                             f�     �  $              end somador_v0arch;5��    $                   Y'                    �    $                    \'                     �    $                    ['                     �    $                    Z'                     �    $                
   Y'             
       5�_�                    �       ����                                                                                                                                                                                                                                                                                                                           #          �          V       f�&     �   �   �       E   #signal c : bit_vector(31 downto 0);       begin           c(0)  <= '0';       c(1)  <= a(0) and b(0);   ;    c(2)  <= (a(1) and b(1)) or (c(1) and (a(1) xor b(1)));   ;    c(3)  <= (a(2) and b(2)) or (c(2) and (a(2) xor b(2)));   ;    c(4)  <= (a(3) and b(3)) or (c(3) and (a(3) xor b(3)));   ;    c(5)  <= (a(4) and b(4)) or (c(4) and (a(4) xor b(4)));   ;    c(6)  <= (a(5) and b(5)) or (c(5) and (a(5) xor b(5)));   ;    c(7)  <= (a(6) and b(6)) or (c(6) and (a(6) xor b(6)));   ;    c(8)  <= (a(7) and b(7)) or (c(7) and (a(7) xor b(7)));   ;    c(9)  <= (a(8) and b(8)) or (c(8) and (a(8) xor b(8)));   ;    c(10) <= (a(9) and b(9)) or (c(9) and (a(9) xor b(9)));   @    c(11) <= (a(10) and b(10)) or (c(10) and (a(10) xor b(10)));   @    c(12) <= (a(11) and b(11)) or (c(11) and (a(11) xor b(11)));   @    c(13) <= (a(12) and b(12)) or (c(12) and (a(12) xor b(12)));   @    c(14) <= (a(13) and b(13)) or (c(13) and (a(13) xor b(13)));   @    c(15) <= (a(14) and b(14)) or (c(14) and (a(14) xor b(14)));   @    c(16) <= (a(15) and b(15)) or (c(15) and (a(15) xor b(15)));   @    c(17) <= (a(16) and b(16)) or (c(16) and (a(16) xor b(16)));   @    c(18) <= (a(17) and b(17)) or (c(17) and (a(17) xor b(17)));   @    c(19) <= (a(18) and b(18)) or (c(18) and (a(18) xor b(18)));   @    c(20) <= (a(19) and b(19)) or (c(19) and (a(19) xor b(19)));   @    c(21) <= (a(20) and b(20)) or (c(20) and (a(20) xor b(20)));   @    c(22) <= (a(21) and b(21)) or (c(21) and (a(21) xor b(21)));   @    c(23) <= (a(22) and b(22)) or (c(22) and (a(22) xor b(22)));   @    c(24) <= (a(23) and b(23)) or (c(23) and (a(23) xor b(23)));   @    c(25) <= (a(24) and b(24)) or (c(24) and (a(24) xor b(24)));   @    c(26) <= (a(25) and b(25)) or (c(25) and (a(25) xor b(25)));   @    c(27) <= (a(26) and b(26)) or (c(26) and (a(26) xor b(26)));   @    c(28) <= (a(27) and b(27)) or (c(27) and (a(27) xor b(27)));   @    c(29) <= (a(28) and b(28)) or (c(28) and (a(28) xor b(28)));   @    c(30) <= (a(29) and b(29)) or (c(29) and (a(29) xor b(29)));   @    c(31) <= (a(30) and b(30)) or (c(30) and (a(30) xor b(30)));             soma(0)  <= a(0) xor b(0);   '    soma(1)  <= a(1) xor b(1) xor c(1);   '    soma(2)  <= a(2) xor b(2) xor c(2);   '    soma(3)  <= a(3) xor b(3) xor c(3);   '    soma(4)  <= a(4) xor b(4) xor c(4);   '    soma(5)  <= a(5) xor b(5) xor c(5);   '    soma(6)  <= a(6) xor b(6) xor c(6);   '    soma(7)  <= a(7) xor b(7) xor c(7);   '    soma(8)  <= a(8) xor b(8) xor c(8);   '    soma(9)  <= a(9) xor b(9) xor c(9);   *    soma(10) <= a(10) xor b(10) xor c(10);   *    soma(11) <= a(11) xor b(11) xor c(11);   *    soma(12) <= a(12) xor b(12) xor c(12);   *    soma(13) <= a(13) xor b(13) xor c(13);   *    soma(14) <= a(14) xor b(14) xor c(14);   *    soma(15) <= a(15) xor b(15) xor c(15);   *    soma(16) <= a(16) xor b(16) xor c(16);   *    soma(17) <= a(17) xor b(17) xor c(17);   *    soma(18) <= a(18) xor b(18) xor c(18);   *    soma(19) <= a(19) xor b(19) xor c(19);   *    soma(20) <= a(20) xor b(20) xor c(20);   *    soma(21) <= a(21) xor b(21) xor c(21);   *    soma(22) <= a(22) xor b(22) xor c(22);   *    soma(23) <= a(23) xor b(23) xor c(23);   *    soma(24) <= a(24) xor b(24) xor c(24);   *    soma(25) <= a(25) xor b(25) xor c(25);   *    soma(26) <= a(26) xor b(26) xor c(26);   *    soma(27) <= a(27) xor b(27) xor c(27);   *    soma(28) <= a(28) xor b(28) xor c(28);   *    soma(29) <= a(29) xor b(29) xor c(29);   *    soma(30) <= a(30) xor b(30) xor c(30);   *    soma(31) <= a(31) xor b(31) xor c(31);5��    �       E               I                    5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�(     �   �   �   �      ,architecture somador_v0arch of somador_v0 is5��    �                 
   )             
       5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�+     �   �   �   �      (architecture behavioral of somador_v0 is5��    �          
       	   7      
       	       5�_�                    �   #    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�?     �   �   �   �          �   �   �   �    �   �   �   �    5��    �                      D                     �    �                      D                     �    �                      D                     �    �                      D                    5�_�      !               �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�B    �   �   �           5��    �                      Y                     5�_�       "           !   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�w     �   �   �   �      end somador_v0;5��    �          
       	         
       	       5�_�   !   #           "   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�{     �   �   �   �      entity somador_v0 is5��    �          
       	   �      
       	       5�_�   "   $           #   �   C    ����                                                                                                                                                                                                                                                                                                                            �   C       �   C          C    f��     �   �   �   �      `        inst7: somador_v0 port map (a => b_out, b => x"bb67ae85",  soma =>  haso(63 downto 32));   `        inst8: somador_v0 port map (a => c_out, b => x"3c6ef372",  soma =>  haso(95 downto 64));   a        inst9: somador_v0 port map (a => d_out, b => x"a54ff53a",  soma =>  haso(127 downto 96));�   �   �   �      _        inst6: somador_v0 port map (a => a_out, b => x"6a09e667",  soma =>  haso(31 downto 0));5��    �   C                  �                     �    �   C                                       �    �   C                  g                     �    �   C                  �                     5�_�   #   %           $   �   E    ����                                                                                                                                                                                                                                                                                                                            �   E       �   G          G    f��     �   �   �   �      `        inst6: somador_v0 port map (a => a_out, b => x"6a09e667",   soma =>  haso(31 downto 0));   a        inst7: somador_v0 port map (a => b_out, b => x"bb67ae85",   soma =>  haso(63 downto 32));   a        inst8: somador_v0 port map (a => c_out, b => x"3c6ef372",   soma =>  haso(95 downto 64));   b        inst9: somador_v0 port map (a => d_out, b => x"a54ff53a",   soma =>  haso(127 downto 96));   b        inst10: somador_v0 port map (a => e_out, b => x"510e527f",  soma => haso(159 downto 128));   b        inst11: somador_v0 port map (a => f_out, b => x"9b05688c",  soma => haso(191 downto 160));   b        inst12: somador_v0 port map (a => g_out, b => x"1f83d9ab",  soma => haso(223 downto 192));   b        inst13: somador_v0 port map (a => h_out, b => x"5be0cd19",  soma => haso(255 downto 224));5��    �   E                  �                     �    �   E                                       �    �   E                  c                     �    �   E                  �                     �    �   E                  "                     �    �   E                  �                     �    �   E                  �                     �    �   E                  B                     5�_�   $   &           %   )       ����                                                                                                                                                                                                                                                                                                                            �   E       �   G          G    f��     �   (   *   �      '        q: _out bit_vector(31 downto 0)5��    (                     :                     5�_�   %   '           &   �   8    ����                                                                                                                                                                                                                                                                                                                            �   E       �   G          G    f��     �   �   �   �      H        	sum: somador_v0 port map(a => waux, b => kaux, soma => kpwaux);5��    �   8                 �                    5�_�   &   (           '   "       ����                                                                                                                                                                                                                                                                                                                            �   E       �   G          G    f��    �   !   #   �      '        q: _out bit_vector(31 downto 0)5��    !                     �                     5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                             f��     �         �      entity multisteps_v0 is5��                         :                      5�_�   (   *           )          ����                                                                                                                                                                                                                                                                                                                                                             f��     �         �      entity multistepsv0 is5��                         :                      5�_�   )   +           *          ����                                                                                                                                                                                                                                                                                                                                                             f��     �         �      entity multisteps0 is5��                         :                      5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                                             f��     �         �      1architecture arqmultisteps_v0 of multisteps_v0 is5��                        �                     �                     
   �              
       �              
          �       
              �                     
   �              
       5�_�   +   -           ,      %    ����                                                                                                                                                                                                                                                                                                                                                             f��     �         �      +architecture behavioral of multisteps_v0 is5��       %                                       5�_�   ,   .           -      %    ����                                                                                                                                                                                                                                                                                                                                                             f��     �         �      *architecture behavioral of multistepsv0 is5��       %                                       5�_�   -   /           .      %    ����                                                                                                                                                                                                                                                                                                                                                             f��     �         �      )architecture behavioral of multisteps0 is5��       %                                       5�_�   .   0           /   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      +        r(i) <= A(i) xor B(i) xor carry(i);5��    �                    z                    5�_�   /   1           0   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      &    soma : out bit_vector(31 downto 0)5��    �                    �                    5�_�   0   2           1   �       ����                                                                                                                                                                                                                                                                                                                                                             f��    �   �   �   �      +    r(31) <= A(31) xor B(31) xor carry(31);5��    �                                        5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                                                             f�     �               �   library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity multisteps is   
    port (           clk, rst: in bit;   +        msgi : in bit_vector(511 downto 0);   ,        haso : out bit_vector(255 downto 0);           done : out bit   );   end entity;       (architecture behavioral of multisteps is       component stepfun is    port (   8  ai,bi,ci,di,ei,fi,gi,hi : in bit_vector (31 downto 0);   "  kpw: in bit_vector(31 downto 0);   7  ao,bo,co,do,eo,fo,go,ho: out bit_vector (31 downto 0)    );    end component;       component somador_v0 is   	    port(   &    a, b : in bit_vector(31 downto 0);   #    s : out bit_vector(31 downto 0)       );   end component;           component sigma0 is    	    port(   &        x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)       );   end component;       component sigma1 is   	    port(   &        x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)       );   end component;       	-- sinais       ?type sinal_array is array (0 to 63) of BIT_VECTOR(31 downto 0);       signal K, W, KPW: sinal_array;   Nsignal ain, bin, cin, din, ein, fin, gin, hin, kpwin: bit_vector(31 downto 0);   Wsignal a_out, b_out, c_out, d_out, e_out, f_out, g_out, h_out: bit_vector(31 downto 0);       	    begin   G    	 -- Inicialização dos valores do sinal com os valores fornecidos       K(0) <= x"428a2f98";       K(1) <= x"71374491";       K(2) <= x"b5c0fbcf";       K(3) <= x"e9b5dba5";       K(4) <= x"3956c25b";       K(5) <= x"59f111f1";       K(6) <= x"923f82a4";       K(7) <= x"ab1c5ed5";       K(8) <= x"d807aa98";       K(9) <= x"12835b01";       K(10) <= x"243185be";       K(11) <= x"550c7dc3";       K(12) <= x"72be5d74";       K(13) <= x"80deb1fe";       K(14) <= x"9bdc06a7";       K(15) <= x"c19bf174";       K(16) <= x"e49b69c1";       K(17) <= x"efbe4786";       K(18) <= x"0fc19dc6";       K(19) <= x"240ca1cc";       K(20) <= x"2de92c6f";       K(21) <= x"4a7484aa";       K(22) <= x"5cb0a9dc";       K(23) <= x"76f988da";       K(24) <= x"983e5152";       K(25) <= x"a831c66d";       K(26) <= x"b00327c8";       K(27) <= x"bf597fc7";       K(28) <= x"c6e00bf3";       K(29) <= x"d5a79147";       K(30) <= x"06ca6351";       K(31) <= x"14292967";       K(32) <= x"27b70a85";       K(33) <= x"2e1b2138";       K(34) <= x"4d2c6dfc";       K(35) <= x"53380d13";       K(36) <= x"650a7354";       K(37) <= x"766a0abb";       K(38) <= x"81c2c92e";       K(39) <= x"92722c85";       K(40) <= x"a2bfe8a1";       K(41) <= x"a81a664b";       K(42) <= x"c24b8b70";       K(43) <= x"c76c51a3";       K(44) <= x"d192e819";       K(45) <= x"d6990624";       K(46) <= x"f40e3585";       K(47) <= x"106aa070";       K(48) <= x"19a4c116";       K(49) <= x"1e376c08";       K(50) <= x"2748774c";       K(51) <= x"34b0bcb5";       K(52) <= x"391c0cb3";       K(53) <= x"4ed8aa4a";       K(54) <= x"5b9cca4f";       K(55) <= x"682e6ff3";       K(56) <= x"748f82ee";       K(57) <= x"78a5636f";       K(58) <= x"84c87814";       K(59) <= x"8cc70208";       K(60) <= x"90befffa";       K(61) <= x"a4506ceb";       K(62) <= x"bef9a3f7";       K(63) <= x"c67178f2";             W(0)  <= msgi(31 downto 0);        W(1)  <= msgi(63 downto 32);        W(2)  <= msgi(95 downto 64);   !    W(3)  <= msgi(127 downto 96);   "    W(4)  <= msgi(159 downto 128);   "    W(5)  <= msgi(191 downto 160);   "    W(6)  <= msgi(223 downto 192);   "    W(7)  <= msgi(255 downto 224);   "    W(8)  <= msgi(287 downto 256);   "    W(9)  <= msgi(319 downto 288);   "    W(10) <= msgi(351 downto 320);   "    W(11) <= msgi(383 downto 352);   "    W(12) <= msgi(415 downto 384);   "    W(13) <= msgi(447 downto 416);   "    W(14) <= msgi(479 downto 448);   "    W(15) <= msgi(511 downto 480);            &    gera_w: for i in 16 to 63 generate   8    	signal y1, y2, y3, y4, y5: bit_vector(31 downto 0);   
    	begin   ,        	inst1: sigma1 port map(W(i-2), y1);   -        	inst2: sigma0 port map(W(i-15), y2);   4        	inst3: somador_v0 port map(y1, W(i-7), y3);   0        	inst4: somador_v0 port map(y3, y2, y4);   5        	inst5: somador_v0 port map(y4, W(i-16), y5);           	W(i) <= y5;       	end generate;              )    gera_kpw: for j in 0 to 63 generate     8    	signal waux, kaux, kpwaux: bit_vector(31 downto 0);           begin           	waux <= W(j);               kaux <= K(j);   E        	sum: somador_v0 port map(a => waux, b => kaux, s => kpwaux);               KPW(j) <= kpwaux;       	end generate;              |        inststep : stepfun port map (ain,bin,cin,din,ein,fin,gin,hin,kpwin,a_out,b_out,c_out,d_out,e_out,f_out,g_out,h_out);              		process(clk)   ,        	variable i : integer range 0 to 64;               begin   '            	if (rising_edge(clk)) then   '                    if (rst = '1') then                           i := 0;   $                        done <= '0';                       end if;       1                    if (rst = '0' and i = 0) then   +                        ain <= x"6a09e667";   +                        bin <= x"bb67ae85";   +                        cin <= x"3c6ef372";   +                        din <= x"a54ff53a";   2                        ein <= x"510e527f";          +                        fin <= x"9b05688c";   +                        gin <= x"1f83d9ab";   +                        hin <= x"5be0cd19";   (                        kpwin <= KPW(0);                       end if;       /                    if (i /= 0 and i < 64) then   %                        ain <= a_out;   %                        bin <= b_out;   %                        cin <= c_out;   %                        din <= d_out;   %                        ein <= e_out;   %                        fin <= f_out;   %                        gin <= g_out;   %                        hin <= h_out;   (                        kpwin <= KPW(i);                       end if;       $                    if (i = 64) then   $                        done <= '1';                       end if;                          2                    if (rst = '0' and i < 64) then                        	i := i + 1;                       end if;                   end if;           end process;               ]        inst6: somador_v0 port map (a => a_out, b => x"6a09e667",   s =>  haso(31 downto 0));   ^        inst7: somador_v0 port map (a => b_out, b => x"bb67ae85",   s =>  haso(63 downto 32));   ^        inst8: somador_v0 port map (a => c_out, b => x"3c6ef372",   s =>  haso(95 downto 64));   _        inst9: somador_v0 port map (a => d_out, b => x"a54ff53a",   s =>  haso(127 downto 96));   _        inst10: somador_v0 port map (a => e_out, b => x"510e527f",  s => haso(159 downto 128));   _        inst11: somador_v0 port map (a => f_out, b => x"9b05688c",  s => haso(191 downto 160));   _        inst12: somador_v0 port map (a => g_out, b => x"1f83d9ab",  s => haso(223 downto 192));   _        inst13: somador_v0 port map (a => h_out, b => x"5be0cd19",  s => haso(255 downto 224));              end architecture;       --somador_v0       entity somador32 is   port(   &    a, b : in bit_vector(31 downto 0);   #    s : out bit_vector(31 downto 0)       );   end somador32;       'architecture behavioral of somador32 is   +    signal carry : bit_vector(31 downto 0);   begin   "    sum: for i in 0 to 30 generate   +        s(i) <= A(i) xor B(i) xor carry(i);   T        carry(i+1) <= (A(i) and B(i)) or (A(i) and carry(i)) or (B(i) and carry(i));       end generate;       +    s(31) <= A(31) xor B(31) xor carry(31);         end behavioral;5�5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                                                       f�     �         �      8  ai,bi,ci,di,ei,fi,gi,hi : in bit_vector (31 downto 0);   "  kpw: in bit_vector(31 downto 0);   7  ao,bo,co,do,eo,fo,go,ho: out bit_vector (31 downto 0)    );�         �       port (5��                         #                     �                         .                     �                         j                     �                         �                     �                         �                     5�_�   3   5           4           ����                                                                                                                                                                                                                                                                                                                                                       f�"     �         �       end component;5��                          �                     5�_�   4   6           5           ����                                                                                                                                                                                                                                                                                                                                       +                   f�)     �      ,   �      
    port (   ;     ai,bi,ci,di,ei,fi,gi,hi : in bit_vector (31 downto 0);   %     kpw: in bit_vector(31 downto 0);   :     ao,bo,co,do,eo,fo,go,ho: out bit_vector (31 downto 0)       );   end component;       component somador_v0 is   	    port(   &    a, b : in bit_vector(31 downto 0);   #    s : out bit_vector(31 downto 0)       );   end component;           component sigma0 is    	    port(   &        x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)       );   end component;       component sigma1 is   	    port(   &        x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)       );   end component;�         �      component stepfun is5��                                               �                          &                     �                          5                     �                          u                     �                          �                     �                          �                     �                          �                     �                          �                     �                                               �                                               �                          ,                     �                          W                     �                                               �                          �                     �                          �                     �                          �                     �                          �                     �                          �                     �                           �                     �    !                      �                     �    "                      $                     �    #                      /                     �    $                      B                     �    %                      G                     �    &                      _                     �    '                      m                     �    (                      �                     �    )                      �                     �    *                      �                     5�_�   5   7           6   -        ����                                                                                                                                                                                                                                                                                                                            -           3                   f�0     �   -   4   �          ?type sinal_array is array (0 to 63) of BIT_VECTOR(31 downto 0);       signal K, W, KPW: sinal_array;   Nsignal ain, bin, cin, din, ein, fin, gin, hin, kpwin: bit_vector(31 downto 0);   Wsignal a_out, b_out, c_out, d_out, e_out, f_out, g_out, h_out: bit_vector(31 downto 0);�   ,   .   �      	-- sinais5��    ,                      �                     �    -                      �                     �    .                      �                     �    /                      9                     �    0                      >                     �    1                      a                     �    2                      �                     5�_�   6   9           7   /   +    ����                                                                                                                                                                                                                                                                                                                            -           3                   f�5     �   .   0   �      C    type sinal_array is array (0 to 63) of BIT_VECTOR(31 downto 0);5��    .   +       
                 
              �    .   -                  "                     �    .   ,                  !                     �    .   +                                      �    .   5                  *                     �    .   4                  )                     �    .   3                  (                     �    .   2                  '                     �    .   1                  &                     �    .   0                  %                     �    .   /                  $                     �    .   .                  #                     �    .   -                  "                     �    .   ,                  !                     �    .   +              
                 
       �    .   +       
       
          
       
       �    .   +       
                 
              �    .   +              
                 
       5�_�   7   :   8       9   1        ����                                                                                                                                                                                                                                                                                                                            -           3                   f�J     �   �   �          (                        kpwin <= KPW(i);�   �   �          (                        kpwin <= KPW(0);�   �   �                      KPW(j) <= kpwaux;�   0   2   �      "    signal K, W, KPW: sinal_array;5��    0                    O                    �    �                    �                    �    �   !                 	                    �    �   !                 �                    5�_�   9   ;           :   1        ����                                                                                                                                                                                                                                                                                                                            -           3                   f�h     �   �   �                  	waux <= W(j);�   �   �                  	W(i) <= y5;�   �   �          5        	inst5: somador_v0 port map(y4, W(i-16), y5);�   �   �          4        	inst3: somador_v0 port map(y1, W(i-7), y3);�   �   �          -        	inst2: sigma0 port map(W(i-15), y2);�   �   �          ,        	inst1: sigma1 port map(W(i-2), y1);�   �   �          "    W(15) <= msgi(511 downto 480);�   �   �          "    W(14) <= msgi(479 downto 448);�   �   �          "    W(13) <= msgi(447 downto 416);�   �   �          "    W(12) <= msgi(415 downto 384);�   �   �          "    W(11) <= msgi(383 downto 352);�   �   �          "    W(10) <= msgi(351 downto 320);�   �   �          "    W(9)  <= msgi(319 downto 288);�      �          "    W(8)  <= msgi(287 downto 256);�   ~   �          "    W(7)  <= msgi(255 downto 224);�   }             "    W(6)  <= msgi(223 downto 192);�   |   ~          "    W(5)  <= msgi(191 downto 160);�   {   }          "    W(4)  <= msgi(159 downto 128);�   z   |          !    W(3)  <= msgi(127 downto 96);�   y   {               W(2)  <= msgi(95 downto 64);�   x   z               W(1)  <= msgi(63 downto 32);�   w   y              W(0)  <= msgi(31 downto 0);�   0   2   �      &    signal K, W, kpw_vec: sinal_array;5��    0                    L                    �    w                    �                    �    x                                        �    y                    2                    �    z                    W                    �    {                    }                    �    |                    �                    �    }                    �                    �    ~                    �                    �                                            �    �                    @                    �    �                    g                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                                        �    �                    *                    �    �                     �                    �    �                                         �    �   (                 J                    �    �   (                 �                    �    �   	                 �                    �    �                    }                    5�_�   :   <           ;   1        ����                                                                                                                                                                                                                                                                                                                            -           3                   f�z     �   �   �                      kaux <= K(j);�   u   w              K(63) <= x"c67178f2";�   t   v              K(62) <= x"bef9a3f7";�   s   u              K(61) <= x"a4506ceb";�   r   t              K(60) <= x"90befffa";�   q   s              K(59) <= x"8cc70208";�   p   r              K(58) <= x"84c87814";�   o   q              K(57) <= x"78a5636f";�   n   p              K(56) <= x"748f82ee";�   m   o              K(55) <= x"682e6ff3";�   l   n              K(54) <= x"5b9cca4f";�   k   m              K(53) <= x"4ed8aa4a";�   j   l              K(52) <= x"391c0cb3";�   i   k              K(51) <= x"34b0bcb5";�   h   j              K(50) <= x"2748774c";�   g   i              K(49) <= x"1e376c08";�   f   h              K(48) <= x"19a4c116";�   e   g              K(47) <= x"106aa070";�   d   f              K(46) <= x"f40e3585";�   c   e              K(45) <= x"d6990624";�   b   d              K(44) <= x"d192e819";�   a   c              K(43) <= x"c76c51a3";�   `   b              K(42) <= x"c24b8b70";�   _   a              K(41) <= x"a81a664b";�   ^   `              K(40) <= x"a2bfe8a1";�   ]   _              K(39) <= x"92722c85";�   \   ^              K(38) <= x"81c2c92e";�   [   ]              K(37) <= x"766a0abb";�   Z   \              K(36) <= x"650a7354";�   Y   [              K(35) <= x"53380d13";�   X   Z              K(34) <= x"4d2c6dfc";�   W   Y              K(33) <= x"2e1b2138";�   V   X              K(32) <= x"27b70a85";�   U   W              K(31) <= x"14292967";�   T   V              K(30) <= x"06ca6351";�   S   U              K(29) <= x"d5a79147";�   R   T              K(28) <= x"c6e00bf3";�   Q   S              K(27) <= x"bf597fc7";�   P   R              K(26) <= x"b00327c8";�   O   Q              K(25) <= x"a831c66d";�   N   P              K(24) <= x"983e5152";�   M   O              K(23) <= x"76f988da";�   L   N              K(22) <= x"5cb0a9dc";�   K   M              K(21) <= x"4a7484aa";�   J   L              K(20) <= x"2de92c6f";�   I   K              K(19) <= x"240ca1cc";�   H   J              K(18) <= x"0fc19dc6";�   G   I              K(17) <= x"efbe4786";�   F   H              K(16) <= x"e49b69c1";�   E   G              K(15) <= x"c19bf174";�   D   F              K(14) <= x"9bdc06a7";�   C   E              K(13) <= x"80deb1fe";�   B   D              K(12) <= x"72be5d74";�   A   C              K(11) <= x"550c7dc3";�   @   B              K(10) <= x"243185be";�   ?   A              K(9) <= x"12835b01";�   >   @              K(8) <= x"d807aa98";�   =   ?              K(7) <= x"ab1c5ed5";�   <   >              K(6) <= x"923f82a4";�   ;   =              K(5) <= x"59f111f1";�   :   <              K(4) <= x"3956c25b";�   9   ;              K(3) <= x"e9b5dba5";�   8   :              K(2) <= x"b5c0fbcf";�   7   9              K(1) <= x"71374491";�   6   8              K(0) <= x"428a2f98";�   0   2   �      *    signal K, w_vec, kpw_vec: sinal_array;5��    0                    I                    �    6                    u                    �    7                    �                    �    8                    �                    �    9                    �                    �    :                    �                    �    ;                                        �    <                    /                    �    =                    N                    �    >                    m                    �    ?                    �                    �    @                    �                    �    A                    �                    �    B                    �                    �    C                                        �    D                    +                    �    E                    K                    �    F                    k                    �    G                    �                    �    H                    �                    �    I                    �                    �    J                    �                    �    K                                        �    L                    +                    �    M                    K                    �    N                    k                    �    O                    �                    �    P                    �                    �    Q                    �                    �    R                    �                    �    S                    	                    �    T                    +	                    �    U                    K	                    �    V                    k	                    �    W                    �	                    �    X                    �	                    �    Y                    �	                    �    Z                    �	                    �    [                    
                    �    \                    +
                    �    ]                    K
                    �    ^                    k
                    �    _                    �
                    �    `                    �
                    �    a                    �
                    �    b                    �
                    �    c                                        �    d                    +                    �    e                    K                    �    f                    k                    �    g                    �                    �    h                    �                    �    i                    �                    �    j                    �                    �    k                                        �    l                    +                    �    m                    K                    �    n                    k                    �    o                    �                    �    p                    �                    �    q                    �                    �    r                    �                    �    s                                        �    t                    +                    �    u                    K                    �    �                    !                    5�_�   ;   >           <   �        ����                                                                                                                                                                                                                                                                                                                            -           3                   f��     �   �   �          !            kpw_vec(j) <= kpwaux;�   �   �          E        	sum: somador_v0 port map(a => waux, b => kaux, s => kpwaux);�   �   �                      kaux <= k_const(j);�   �   �                  	waux <= w_vec(j);�   �   �   �      8    	signal waux, kaux, kpwaux: bit_vector(31 downto 0);5��    �                    �                    �    �                    �                    �    �                    �                    �    �   
                 �                    �    �                                        �    �   (                 Z                    �    �   4                 f                    �    �   B                 t                    �    �                    �                    5�_�   <   ?   =       >   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      _        inst10: somador_v0 port map (a => e_out, b => x"510e527f",  s => haso(159 downto 128));   _        inst11: somador_v0 port map (a => f_out, b => x"9b05688c",  s => haso(191 downto 160));   _        inst12: somador_v0 port map (a => g_out, b => x"1f83d9ab",  s => haso(223 downto 192));   _        inst13: somador_v0 port map (a => h_out, b => x"5be0cd19",  s => haso(255 downto 224));5��    �                     x                     �    �                     �                     �    �                     6                     �    �                     �                     5�_�   >   A           ?   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      X        : somador_v0 port map (a => a_out, b => x"6a09e667",   s =>  haso(31 downto 0));�   �   �   �      ]        inst6: somador_v0 port map (a => a_out, b => x"6a09e667",   s =>  haso(31 downto 0));   ^        inst7: somador_v0 port map (a => b_out, b => x"bb67ae85",   s =>  haso(63 downto 32));   ^        inst8: somador_v0 port map (a => c_out, b => x"3c6ef372",   s =>  haso(95 downto 64));   _        inst9: somador_v0 port map (a => d_out, b => x"a54ff53a",   s =>  haso(127 downto 96));   ^        inst1: somador_v0 port map (a => e_out, b => x"510e527f",  s => haso(159 downto 128));   ^        inst1: somador_v0 port map (a => f_out, b => x"9b05688c",  s => haso(191 downto 160));   ^        inst1: somador_v0 port map (a => g_out, b => x"1f83d9ab",  s => haso(223 downto 192));   ^        inst1: somador_v0 port map (a => h_out, b => x"5be0cd19",  s => haso(255 downto 224));5��    �                     �                     �    �                     P                     �    �                     �                     �    �                                          �    �                     _                     �    �                     �                     �    �                                          �    �                     m                     �    �                     �                     �    �                     U                     �    �                     �                     �    �                                          �    �                     s                     �    �                     �                     �    �                     1                     �    �                     �                     5�_�   ?   B   @       A   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      ^        get_a: somador_v0 port map (a => b_out, b => x"bb67ae85",   s =>  haso(63 downto 32));   ^        get_a: somador_v0 port map (a => c_out, b => x"3c6ef372",   s =>  haso(95 downto 64));   _        get_a: somador_v0 port map (a => d_out, b => x"a54ff53a",   s =>  haso(127 downto 96));   ^        get_a: somador_v0 port map (a => e_out, b => x"510e527f",  s => haso(159 downto 128));   ^        get_a: somador_v0 port map (a => f_out, b => x"9b05688c",  s => haso(191 downto 160));   ^        get_a: somador_v0 port map (a => g_out, b => x"1f83d9ab",  s => haso(223 downto 192));   ^        get_a: somador_v0 port map (a => h_out, b => x"5be0cd19",  s => haso(255 downto 224));�   �   �   �      ]        get_a: somador_v0 port map (a => a_out, b => x"6a09e667",   s =>  haso(31 downto 0));5��    �                     �                     �    �                     ]                     �    �                     �                     �    �                     !                     �    �                     �                     �    �                     �                     �    �                     H                     �    �                     �                     5�_�   A   C           B   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      a        get_aout: somador_v0 port map (a => b_out, b => x"bb67ae85",   s =>  haso(63 downto 32));5��    �                    \                    5�_�   B   D           C   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      a        get_aout: somador_v0 port map (a => c_out, b => x"3c6ef372",   s =>  haso(95 downto 64));5��    �                    �                    5�_�   C   E           D   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      b        get_aout: somador_v0 port map (a => d_out, b => x"a54ff53a",   s =>  haso(127 downto 96));5��    �                                         5�_�   D   F           E   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      a        get_aout: somador_v0 port map (a => e_out, b => x"510e527f",  s => haso(159 downto 128));5��    �                    �                    5�_�   E   G           F   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      a        get_aout: somador_v0 port map (a => f_out, b => x"9b05688c",  s => haso(191 downto 160));5��    �                    �                    5�_�   F   H           G   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      a        get_aout: somador_v0 port map (a => g_out, b => x"1f83d9ab",  s => haso(223 downto 192));5��    �                    G                    5�_�   G   I           H   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      a        get_aout: somador_v0 port map (a => h_out, b => x"5be0cd19",  s => haso(255 downto 224));5��    �                    �                    5�_�   H   J           I           ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �          "    sum: for i in 0 to 30 generate�   �   �          begin�   �   �          &    a, b : in bit_vector(31 downto 0);�   �   �          ,                        kpwin <= kpw_vec(i);�   �   �          %                        hin <= h_out;�   �   �          %                        gin <= g_out;�   �   �          %                        fin <= f_out;�   �   �          %                        ein <= e_out;�   �   �          %                        din <= d_out;�   �   �          %                        cin <= c_out;�   �   �          %                        bin <= b_out;�   �   �          %                        ain <= a_out;�   �   �          ,                        kpwin <= kpw_vec(0);�   �   �          +                        hin <= x"5be0cd19";�   �   �          +                        gin <= x"1f83d9ab";�   �   �          +                        fin <= x"9b05688c";�   �   �          2                        ein <= x"510e527f";       �   �   �          +                        din <= x"a54ff53a";�   �   �          +                        cin <= x"3c6ef372";�   �   �          +                        bin <= x"bb67ae85";�   �   �          +                        ain <= x"6a09e667";�   �   �          '            	if (rising_edge(clk)) then�   �   �                      begin�   �   �          ,        	variable i : integer range 0 to 64;�   �   �          |        inststep : stepfun port map (ain,bin,cin,din,ein,fin,gin,hin,kpwin,a_out,b_out,c_out,d_out,e_out,f_out,g_out,h_out);�   �   �                  begin�   �   �          )    gera_kpw: for j in 0 to 63 generate  �   �   �          9        	inst5: somador_v0 port map(y4, w_vec(i-16), y5);�   �   �          0        	inst4: somador_v0 port map(y3, y2, y4);�   �   �          8        	inst3: somador_v0 port map(y1, w_vec(i-7), y3);�   �   �          1        	inst2: sigma0 port map(w_vec(i-15), y2);�   �   �          0        	inst1: sigma1 port map(w_vec(i-2), y1);�   �   �          
    	begin�   �   �          &    gera_w: for i in 16 to 63 generate�   5   7          G    	 -- Inicialização dos valores do sinal com os valores fornecidos�   4   6          	    begin�   1   3          R    signal ain, bin, cin, din, ein, fin, gin, hin, kpwin: bit_vector(31 downto 0);�   0   2          0    signal k_const, w_vec, kpw_vec: sinal_array;�   .   0          C    type sinal_array is array (0 to 63) of bit_vector(31 downto 0);�   ,   .              -- sinais�   '   )          *            x: in bit_vector(31 downto 0);�       "          *            x: in bit_vector(31 downto 0);�                *        a, b : in bit_vector(31 downto 0);�                )         kpw: in bit_vector(31 downto 0);�                ?         ai,bi,ci,di,ei,fi,gi,hi : in bit_vector (31 downto 0);�                +        msgi : in bit_vector(511 downto 0);�         �              clk, rst: in bit;5��                        [                     �                        s                     �       #                 Z                    �                        �                    �                        ?                    �                         �                    �    '                    �                    �    ,                    �                    �    .   
                                     �    0   %                 l                    �    1                    �                    �    1                    �                    �    1                    �                    �    1                    �                    �    1   $                 �                    �    1   *                 �                    �    1   0                 �                    �    1   6                 �                    �    1   >                 �                    �    4                    9                    �    5   )                 f                    �    �                                        �    �                    X                    �    �   	                 e                    �    �   	                 �                    �    �   	                 �                    �    �   	                                     �    �   	                 6                    �    �                    �                    �    �                                        �    �                    �                    �    �   '                 �                    �    �   ,                                     �    �   1                 	                    �    �   6                                     �    �   ;                                     �    �   @                                     �    �   E                                     �    �   J                 "                    �    �   Q                 )                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                                        �    �                    =                    �    �                    j                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    '                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                                        �    �                    <                    �    �                    c                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    :                    �    �                    M                    5�_�   I   K           J   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      #    sum: for i _in 0 to 30 generate5��    �                     M                     5�_�   J   L           K          ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �         �              clk, rst: _in bit;5��                         [                      5�_�   K   M           L          ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �         �      ,        msgi : _in bit_vector(511 downto 0);5��                         r                      5�_�   L   N           M      #    ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �         �      @         ai,bi,ci,di,ei,fi,gi,hi : _in bit_vector (31 downto 0);5��       #                  X                     5�_�   M   O           N          ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �         �      *         kpw: _in bit_vector(31 downto 0);5��                         �                     5�_�   N   P           O          ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �         �      +        a, b : _in bit_vector(31 downto 0);5��                         ;                     5�_�   O   Q           P   !       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �       "   �      +            x: _in bit_vector(31 downto 0);5��                          �                     5�_�   P   R           Q   (       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   '   )   �      +            x: _in bit_vector(31 downto 0);5��    '                     |                     5�_�   Q   S           R   5       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   4   6   �      
    beg_in5��    4                     2                     5�_�   R   U           S   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      '    gera_w: for i _in 16 to 63 generate5��    �                     �                     5�_�   S   V   T       U   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f�     �   �   �   �          	beg_in5��    �                     O                     5�_�   U   W           V   �   	    ����                                                                                                                                                                                                                                                                                                                            �   	       �   	              f�
     �   �   �   �      1        	_inst1: sigma1 port map(w_vec(i-2), y1);   2        	_inst2: sigma0 port map(w_vec(i-15), y2);   9        	_inst3: somador_v0 port map(y1, w_vec(i-7), y3);   1        	_inst4: somador_v0 port map(y3, y2, y4);   :        	_inst5: somador_v0 port map(y4, w_vec(i-16), y5);5��    �   	                  [                     �    �   	                  �                     �    �   	                  �                     �    �   	                  �                     �    �   	                  (                     5�_�   V   X           W   �   	    ����                                                                                                                                                                                                                                                                                                                            �   	       �                 f�     �   �   �   �      ,        	1: sigma1 port map(w_vec(i-2), y1);�   �   �   �      0        	inst1: sigma1 port map(w_vec(i-2), y1);   1        	inst2: sigma0 port map(w_vec(i-15), y2);   8        	inst3: somador_v0 port map(y1, w_vec(i-7), y3);   0        	inst4: somador_v0 port map(y3, y2, y4);   9        	inst5: somador_v0 port map(y4, w_vec(i-16), y5);5��    �   	                  [                     �    �   	                  �                     �    �   	                  �                     �    �   	                  �                     �    �   	                                       �    �   	                  [                     �    �   	                  �                     �    �   	                  �                     �    �   	                  �                     �    �   	                  (                     5�_�   W   Y           X   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�     �   �   �                  	w_vec(i) <= y5;�   �   �          9        	make5: somador_v0 port map(y4, w_vec(i-16), y5);�   �   �          0        	make4: somador_v0 port map(y3, y2, y4);�   �   �          8        	make3: somador_v0 port map(y1, w_vec(i-7), y3);�   �   �          1        	make2: sigma0 port map(w_vec(i-15), y2);�   �   �          0        	make1: sigma1 port map(w_vec(i-2), y1);�   �   �   �      8    	signal y1, y2, y3, y4, y5: bit_vector(31 downto 0);5��    �                                        �    �                                        �    �                    $                    �    �                    )                    �    �                     .                    �    �   ,                 �                    �    �   -                 �                    �    �   $                 �                    �    �   5                 �                    �    �   $                                     �    �   )                                      �    �   .                 %                    �    �   $                 O                    �    �   6                 a                    �    �                    |                    5�_�   X   Z           Y   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�      �   �   �   �              beg_in5��    �                                          5�_�   Y   [           Z   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�#     �   �   �   �      *    gera_kpw: for j _in 0 to 63 generate  5��    �                     �                     5�_�   Z   \           [   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�)     �   �   �   �      �        _inststep : stepfun port map (a_in,b_in,c_in,d_in,e_in,f_in,g_in,h_in,kpw_in,a_out,b_out,c_out,d_out,e_out,f_out,g_out,h_out);5��    �                     �                     5�_�   [   ]           \   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�*     �   �   �   �      �        inststep : stepfun port map (a_in,b_in,c_in,d_in,e_in,f_in,g_in,h_in,kpw_in,a_out,b_out,c_out,d_out,e_out,f_out,g_out,h_out);5��    �                     �                     5�_�   \   ^           ]   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�*     �   �   �   �      �        nststep : stepfun port map (a_in,b_in,c_in,d_in,e_in,f_in,g_in,h_in,kpw_in,a_out,b_out,c_out,d_out,e_out,f_out,g_out,h_out);5��    �                     �                     5�_�   ]   _           ^   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�+     �   �   �   �      �        ststep : stepfun port map (a_in,b_in,c_in,d_in,e_in,f_in,g_in,h_in,kpw_in,a_out,b_out,c_out,d_out,e_out,f_out,g_out,h_out);5��    �                     �                     5�_�   ^   `           _   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�+     �   �   �   �      �        tstep : stepfun port map (a_in,b_in,c_in,d_in,e_in,f_in,g_in,h_in,kpw_in,a_out,b_out,c_out,d_out,e_out,f_out,g_out,h_out);5��    �                     �                     5�_�   _   a           `   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�,     �   �   �   �      �        step : stepfun port map (a_in,b_in,c_in,d_in,e_in,f_in,g_in,h_in,kpw_in,a_out,b_out,c_out,d_out,e_out,f_out,g_out,h_out);5��    �                     �                     5�_�   `   b           a   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�1     �   �   �   �                  beg_in5��    �                     �                     5�_�   a   c           b   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�2     �   �   �   �      -        	variable i : _integer range 0 to 64;5��    �                     �                     5�_�   b   d           c   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�6     �   �   �   �      '    a, b : _in bit_vector(31 downto 0);5��    �                     �                     5�_�   c   e           d   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�8     �   �   �   �      beg_in5��    �                     5                     5�_�   d   f           e   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�;   	 �   �   �   �      (            	if (ris_ing_edge(clk)) then5��    �                     �                     5�_�   e   g           f           ����                                                                                                                                                                                                                                                                                                                                       �           V        f��     �              �   library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity multisteps is   
    port (           clk, rst: in bit;   +        msgi : in bit_vector(511 downto 0);   ,        haso : out bit_vector(255 downto 0);           done : out bit   );   end entity;       (architecture behavioral of multisteps is           component stepfun is           port (   ?         ai,bi,ci,di,ei,fi,gi,hi : in bit_vector (31 downto 0);   )         kpw: in bit_vector(31 downto 0);   >         ao,bo,co,do,eo,fo,go,ho: out bit_vector (31 downto 0)   
        );       end component;               component somador_v0 is           port(   *        a, b : in bit_vector(31 downto 0);   '        s : out bit_vector(31 downto 0)   
        );       end component;                     component sigma0 is            port(   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;              component sigma1 is           port(   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           -- s_inais          D    type s_inal_array is array (0 to 63) of bit_vector(31 downto 0);          1    signal k_const, w_vec, kpw_vec: s_inal_array;   [    signal a_in, b_in, c_in, d_in, e_in, f_in, g_in, h_in, kpw_in: bit_vector(31 downto 0);   [    signal a_out, b_out, c_out, d_out, e_out, f_out, g_out, h_out: bit_vector(31 downto 0);       	    begin   H    	 -- Inicialização dos valores do s_inal com os valores fornecidos       k_const(0) <= x"428a2f98";       k_const(1) <= x"71374491";       k_const(2) <= x"b5c0fbcf";       k_const(3) <= x"e9b5dba5";       k_const(4) <= x"3956c25b";       k_const(5) <= x"59f111f1";       k_const(6) <= x"923f82a4";       k_const(7) <= x"ab1c5ed5";       k_const(8) <= x"d807aa98";       k_const(9) <= x"12835b01";       k_const(10) <= x"243185be";       k_const(11) <= x"550c7dc3";       k_const(12) <= x"72be5d74";       k_const(13) <= x"80deb1fe";       k_const(14) <= x"9bdc06a7";       k_const(15) <= x"c19bf174";       k_const(16) <= x"e49b69c1";       k_const(17) <= x"efbe4786";       k_const(18) <= x"0fc19dc6";       k_const(19) <= x"240ca1cc";       k_const(20) <= x"2de92c6f";       k_const(21) <= x"4a7484aa";       k_const(22) <= x"5cb0a9dc";       k_const(23) <= x"76f988da";       k_const(24) <= x"983e5152";       k_const(25) <= x"a831c66d";       k_const(26) <= x"b00327c8";       k_const(27) <= x"bf597fc7";       k_const(28) <= x"c6e00bf3";       k_const(29) <= x"d5a79147";       k_const(30) <= x"06ca6351";       k_const(31) <= x"14292967";       k_const(32) <= x"27b70a85";       k_const(33) <= x"2e1b2138";       k_const(34) <= x"4d2c6dfc";       k_const(35) <= x"53380d13";       k_const(36) <= x"650a7354";       k_const(37) <= x"766a0abb";       k_const(38) <= x"81c2c92e";       k_const(39) <= x"92722c85";       k_const(40) <= x"a2bfe8a1";       k_const(41) <= x"a81a664b";       k_const(42) <= x"c24b8b70";       k_const(43) <= x"c76c51a3";       k_const(44) <= x"d192e819";       k_const(45) <= x"d6990624";       k_const(46) <= x"f40e3585";       k_const(47) <= x"106aa070";       k_const(48) <= x"19a4c116";       k_const(49) <= x"1e376c08";       k_const(50) <= x"2748774c";       k_const(51) <= x"34b0bcb5";       k_const(52) <= x"391c0cb3";       k_const(53) <= x"4ed8aa4a";       k_const(54) <= x"5b9cca4f";       k_const(55) <= x"682e6ff3";       k_const(56) <= x"748f82ee";       k_const(57) <= x"78a5636f";       k_const(58) <= x"84c87814";       k_const(59) <= x"8cc70208";       k_const(60) <= x"90befffa";       k_const(61) <= x"a4506ceb";       k_const(62) <= x"bef9a3f7";       k_const(63) <= x"c67178f2";         #    w_vec(0)  <= msgi(31 downto 0);   $    w_vec(1)  <= msgi(63 downto 32);   $    w_vec(2)  <= msgi(95 downto 64);   %    w_vec(3)  <= msgi(127 downto 96);   &    w_vec(4)  <= msgi(159 downto 128);   &    w_vec(5)  <= msgi(191 downto 160);   &    w_vec(6)  <= msgi(223 downto 192);   &    w_vec(7)  <= msgi(255 downto 224);   &    w_vec(8)  <= msgi(287 downto 256);   &    w_vec(9)  <= msgi(319 downto 288);   &    w_vec(10) <= msgi(351 downto 320);   &    w_vec(11) <= msgi(383 downto 352);   &    w_vec(12) <= msgi(415 downto 384);   &    w_vec(13) <= msgi(447 downto 416);   &    w_vec(14) <= msgi(479 downto 448);   &    w_vec(15) <= msgi(511 downto 480);            &    gera_w: for i in 16 to 63 generate   =    	signal op1, op2, op3, op4, op5: bit_vector(31 downto 0);   
    	begin   1        	make1: sigma1 port map(w_vec(i-2), op1);   2        	make2: sigma0 port map(w_vec(i-15), op2);   :        	make3: somador_v0 port map(op1, w_vec(i-7), op3);   3        	make4: somador_v0 port map(op3, op2, op4);   ;        	make5: somador_v0 port map(op4, w_vec(i-16), op5);           	w_vec(i) <= op5;       	end generate;              )    gera_kpw: for j in 0 to 63 generate     ;    	signal w_aux, k_aux, kpw_aux: bit_vector(31 downto 0);           begin           	w_aux <= w_vec(j);                k_aux <= k_const(j);   H        	sum: somador_v0 port map(a => w_aux, b => k_aux, s => kpw_aux);   "            kpw_vec(j) <= kpw_aux;       	end generate;              �        make_step : stepfun port map (a_in,b_in,c_in,d_in,e_in,f_in,g_in,h_in,kpw_in,a_out,b_out,c_out,d_out,e_out,f_out,g_out,h_out);              		process(clk)   ,        	variable i : integer range 0 to 64;               begin   '            	if (rising_edge(clk)) then   '                    if (rst = '1') then                           i := 0;   $                        done <= '0';                       end if;       1                    if (rst = '0' and i = 0) then   ,                        a_in <= x"6a09e667";   ,                        b_in <= x"bb67ae85";   ,                        c_in <= x"3c6ef372";   ,                        d_in <= x"a54ff53a";   3                        e_in <= x"510e527f";          ,                        f_in <= x"9b05688c";   ,                        g_in <= x"1f83d9ab";   ,                        h_in <= x"5be0cd19";   -                        kpw_in <= kpw_vec(0);                       end if;       /                    if (i /= 0 and i < 64) then   &                        a_in <= a_out;   &                        b_in <= b_out;   &                        c_in <= c_out;   &                        d_in <= d_out;   &                        e_in <= e_out;   &                        f_in <= f_out;   &                        g_in <= g_out;   &                        h_in <= h_out;   -                        kpw_in <= kpw_vec(i);                       end if;       $                    if (i = 64) then   $                        done <= '1';                       end if;                          2                    if (rst = '0' and i < 64) then                        	i := i + 1;                       end if;                   end if;           end process;               `        get_aout: somador_v0 port map (a => a_out, b => x"6a09e667",   s =>  haso(31 downto 0));   a        get_bout: somador_v0 port map (a => b_out, b => x"bb67ae85",   s =>  haso(63 downto 32));   a        get_cout: somador_v0 port map (a => c_out, b => x"3c6ef372",   s =>  haso(95 downto 64));   b        get_dout: somador_v0 port map (a => d_out, b => x"a54ff53a",   s =>  haso(127 downto 96));   a        get_eout: somador_v0 port map (a => e_out, b => x"510e527f",  s => haso(159 downto 128));   a        get_fout: somador_v0 port map (a => f_out, b => x"9b05688c",  s => haso(191 downto 160));   a        get_gout: somador_v0 port map (a => g_out, b => x"1f83d9ab",  s => haso(223 downto 192));   a        get_hout: somador_v0 port map (a => h_out, b => x"5be0cd19",  s => haso(255 downto 224));              end architecture;       --somador_v0       entity somador32 is   port(   &    a, b : in bit_vector(31 downto 0);   #    s : out bit_vector(31 downto 0)       );   end somador32;       'architecture behavioral of somador32 is   +    signal carry : bit_vector(31 downto 0);   begin   "    sum: for i in 0 to 30 generate   +        s(i) <= A(i) xor B(i) xor carry(i);   T        carry(i+1) <= (A(i) and B(i)) or (A(i) and carry(i)) or (B(i) and carry(i));       end generate;       +    s(31) <= A(31) xor B(31) xor carry(31);         end behavioral;5��            �                      .             5�_�   f   h           g           ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �                  gera_w: for i i�   �            �                   �               5��                    �                      �      �    �              a       �              )      5�_�   g   i           h   �        ����                                                                                                                                                                                                                                                                                                                                                  V        f��    �   �   �           5��    �                      "                     5�_�   h   j           i   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        f��     �   �   �          entity somador32 is   port(   &    a, b : in bit_vector(31 downto 0);   #    s : out bit_vector(31 downto 0)       );   end somador32;       'architecture behavioral of somador32 is   +    signal carry : bit_vector(31 downto 0);   begin   "    sum: for i in 0 to 30 generate   +        s(i) <= A(i) xor B(i) xor carry(i);   T        carry(i+1) <= (A(i) and B(i)) or (A(i) and carry(i)) or (B(i) and carry(i));       end generate;       +    s(31) <= A(31) xor B(31) xor carry(31);         end behavioral;5��    �                      T      �              5�_�   i   k           j          ����                                                                                                                                                                                                                                                                                                                            �           �           V        f��    �         �      entity multisteps is5��                         :                      5�_�   j   l           k      %    ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�    �         �      (architecture behavioral of multisteps is5��       %                                       5�_�   k   m           l   �   &    ����                                                                                                                                                                                                                                                                                                                                                             f�^     �   �   �   �      &    w_vec(15) <= msgi(511 downto 480);5��    �   &                  �                     �    �   )                 �                    �    �   (                  �                     �    �   &                  �                     5�_�   l   n           m   �   &    ����                                                                                                                                                                                                                                                                                                                                                             f�h     �   �   �   �      &    w_vec(15) <= msgi(511 downto 480);5��    �   &                  �                     5�_�   m   p           n   �   &    ����                                                                                                                                                                                                                                                                                                                                                             f�q     �   w   y   �      #    w_vec(0)  <= msgi(31 downto 0);�   x   z   �      $    w_vec(1)  <= msgi(63 downto 32);�   y   {   �      $    w_vec(2)  <= msgi(95 downto 64);�   z   |   �      %    w_vec(3)  <= msgi(127 downto 96);�   {   }   �      &    w_vec(4)  <= msgi(159 downto 128);�   |   ~   �      &    w_vec(5)  <= msgi(191 downto 160);�   }      �      &    w_vec(6)  <= msgi(223 downto 192);�   ~   �   �      &    w_vec(7)  <= msgi(255 downto 224);�      �   �      &    w_vec(8)  <= msgi(287 downto 256);�   �   �   �      &    w_vec(9)  <= msgi(319 downto 288);�   �   �   �      &    w_vec(10) <= msgi(351 downto 320);�   �   �   �      &    w_vec(11) <= msgi(383 downto 352);�   �   �   �      &    w_vec(12) <= msgi(415 downto 384);�   �   �   �      &    w_vec(13) <= msgi(447 downto 416);�   �   �   �      &    w_vec(14) <= msgi(479 downto 448);5��    �   &                  �                     �    �   &                  �                     �    �   &                  o                     �    �   &                  H                     �    �   &                  !                     �    �   &                  �                     �       &                  �                     �    ~   &                  �                     �    }   &                  �                     �    |   &                  ^                     �    {   &                  7                     �    z   %                                       �    y   $                  �                     �    x   $                  �                     �    w   #                  �                     5�_�   n   q   o       p   �   +    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �   �   �   �      +    w_vec(14) <= msgi(479 downto 448); -- 05��    �   *                                     5�_�   p   r           q   �   +    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �   �   �   �      +    w_vec(13) <= msgi(447 downto 416); -- 05��    �   *                 �                    5�_�   q   s           r   �   +    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �   �   �   �      +    w_vec(12) <= msgi(415 downto 384); -- 05��    �   *                 �                    5�_�   r   t           s   �   +    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �   �   �   �      +    w_vec(11) <= msgi(383 downto 352); -- 05��    �   *                 �                    �    �   +                  �                     5�_�   s   u           t   �   +    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �   �   �   �      +    w_vec(10) <= msgi(351 downto 320); -- 05��    �   *                 W                    5�_�   t   v           u   �   *    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �   �   �   �      +    w_vec(9)  <= msgi(319 downto 288); -- 05��    �   *                 +                    5�_�   u   w           v   �   *    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �      �   �      +    w_vec(8)  <= msgi(287 downto 256); -- 05��       *                 �                    5�_�   v   x           w      *    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �   ~   �   �      +    w_vec(7)  <= msgi(255 downto 224); -- 05��    ~   *                 �                    5�_�   w   y           x   ~   *    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �   }      �      +    w_vec(6)  <= msgi(223 downto 192); -- 05��    }   *                 �                    5�_�   x   z           y   }   *    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �   |   ~   �      +    w_vec(5)  <= msgi(191 downto 160); -- 05��    |   *                 {                    5�_�   y   {           z   }   +    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �   |   ~   �      +    w_vec(5)  <= msgi(191 downto 160); -- 15��    |   +                  |                     5�_�   z   |           {   |   +    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �   {   }   �      +    w_vec(4)  <= msgi(159 downto 128); -- 05��    {   *                 O                    5�_�   {   }           |   {   *    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �   z   |   �      *    w_vec(3)  <= msgi(127 downto 96); -- 05��    z   )                 #                    5�_�   |   ~           }   z   )    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �   y   {   �      )    w_vec(2)  <= msgi(95 downto 64); -- 05��    y   (                 �                    5�_�   }              ~   y   )    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��     �   x   z   �      )    w_vec(1)  <= msgi(63 downto 32); -- 05��    x   (                 �                    5�_�   ~                  x   (    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f��    �   w   y   �      (    w_vec(0)  <= msgi(31 downto 0); -- 05��    w   '                 �                    5�_�   n           p   o   x   '    ����                                                                                                                                                                                                                                                                                                                            x   '       �   +       ���    f�}     �   w   �   �      (    w_vec(0)  <= msgi(31 downto 0); -- 1   )    w_vec(1)  <= msgi(63 downto 32); -- 2   )    w_vec(2)  <= msgi(95 downto 64); -- 3   *    w_vec(3)  <= msgi(127 downto 96); -- 4   +    w_vec(4)  <= msgi(159 downto 128); -- 5   +    w_vec(5)  <= msgi(191 downto 160); -- 6   +    w_vec(6)  <= msgi(223 downto 192); -- 7   +    w_vec(7)  <= msgi(255 downto 224); -- 8   +    w_vec(8)  <= msgi(287 downto 256); -- 9   ,    w_vec(9)  <= msgi(319 downto 288); -- 10   ,    w_vec(10) <= msgi(351 downto 320); -- 11   ,    w_vec(11) <= msgi(383 downto 352); -- 12   ,    w_vec(12) <= msgi(415 downto 384); -- 13   ,    w_vec(13) <= msgi(447 downto 416); -- 14   ,    w_vec(14) <= msgi(479 downto 448); -- 155��    w   '                 �                    �    x   (                 �                    �    y   (                 �                    �    z   )                 #                    �    {   *                 O                    �    |   *                 {                    �    }   *                 �                    �    ~   *                 �                    �       *                 �                    �    �   *                 +                    �    �   *                 X                    �    �   *                 �                    �    �   *                 �                    �    �   *                 �                    �    �   *                                     5�_�   S           U   T   �   	    ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      
    	beg_n5��    �   	                  P                     5�_�   ?           A   @   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      `        get_aout: somador_v0 port map (a => a_out, b => x"6a09e667",   s =>  haso(31 downto 0));5��    �                     �                     5�_�   <           >   =   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      ^        inst6 : somador_v0 port map (a => a_out, b => x"6a09e667",   s =>  haso(31 downto 0));�   �   �   �      _        inst7 : somador_v0 port map (a => b_out, b => x"bb67ae85",   s =>  haso(63 downto 32));   _        inst8 : somador_v0 port map (a => c_out, b => x"3c6ef372",   s =>  haso(95 downto 64));   `        inst9 : somador_v0 port map (a => d_out, b => x"a54ff53a",   s =>  haso(127 downto 96));5��    �                     �                     �    �                     [                     �    �                     �                     �    �                                          5�_�   7           9   8   1       ����                                                                                                                                                                                                                                                                                                                            -           3                   f�:     �   0   2   �      "    signal K, W, kpw: sinal_array;5��    0                    O                    5�_�                    �   #    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�8     �   �   �   �    �   �   �   �      1architecture behavioral of somador32somador_v0 is5��    �   $               
   @              
       5�_�   	       
                 ����                                                                                                                                                                                                                                                                                                                            �   G       �   G       V   G    f6�     �        '      component somador_v0 is�   �   �          4        	inst3: somador_v0 port map(y1, W(i-7), y3);�   �   �          0        	inst4: somador_v0 port map(y3, y2, y4);�   �   �          5        	inst5: somador_v0 port map(y4, W(i-16), y5);�   �   �          H        	sum: somador_v0 port map(a => waux, b => kaux, soma => kpwaux);�   �   �          ]        inst6: somador_v0 port map (a => aout, b => x"6a09e667",  soma => haso(31 downto 0));�   �   �          ^        inst7: somador_v0 port map (a => bout, b => x"bb67ae85",  soma => haso(63 downto 32));�   �   �          ^        inst8: somador_v0 port map (a => cout, b => x"3c6ef372",  soma => haso(95 downto 64));�   �   �          _        inst9: somador_v0 port map (a => dout, b => x"a54ff53a",  soma => haso(127 downto 96));�   �   �          a        inst10: somador_v0 port map (a => eout, b => x"510e527f",  soma => haso(159 downto 128));�   �   �          a        inst11: somador_v0 port map (a => fout, b => x"9b05688c",  soma => haso(191 downto 160));�   �   �          a        inst12: somador_v0 port map (a => gout, b => x"1f83d9ab",  soma => haso(223 downto 192));�   �   �          a        inst13: somador_v0 port map (a => hout, b => x"5be0cd19",  soma => haso(255 downto 224));�   �   �          --somador_v0�   �   �          entity somador_v0 is�   �   �          end somador_v0;�   �   �          )architecture somador_v0arch of somador is�  &  (          end somador_v0arch;5��       
              
   �             
       �    �                 
   �             
       �    �                 
   �             
       �    �                 
                
       �    �                 
                
       �    �                 
   �             
       �    �                 
                
       �    �                 
   x             
       �    �                 
   �             
       �    �                 
   8             
       �    �                 
   �             
       �    �                 
   �             
       �    �                 
   ^             
       �    �                 
   �             
       �    �                 
   �             
       �    �                 
   N             
       �    �                 
   h             
       �    &                
   �'             
       5�_�   	              
   �       ����                                                                                                                                                                                                                                                                                                                            �   G       �   G       V   G    f6~     �   �   �  '      entity somadorr is5��    �                     �                     5��