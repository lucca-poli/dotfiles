Vim�UnDo� ��yU�Y.F�	�����W^ ҢU�����   �   A                            serial_o <= not par(0); -- parity bit   �   ,                   fD7   ! _�                             ����                                                                                                                                                                                                                                                                                                                                                             f?#     �                   �               5��                                         �      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f?$     �                  5��                                                  5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f?)     �               5��                          �                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f?)     �                  5��                          �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f?*     �                 end architecture �               architecture rtl of  is�                     �                 arch�                 []5��                          �                     �                          �                     �                          �                     �                          �                     �                         �                     �                         �                    �                         �                    �                         �                    �                         �                    �                        �                     �                          �                      �                        �                     �                         �                     �                         �                     �                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f?-     �             �                 end architecture rtl;�             �             �             �             �             �             �             �             �             �               architecture rtl of tx is5��                        �                    �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                     	   �             	       �                         �                     �              	       
   �      	       
       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f?2     �                architecture Behavioral of tx is5��                        �                    �                         �                     �                         �                     �                         �                     �                     
   �             
       �              
          �      
              �                     
   �             
       5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                v       f?h     �                   �             �                   �             5��                          �                     �                          �                     �                         �                     �                     B   �              =      5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                v       f?m     �                    1.5��                          �                     5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                v       f?n     �                2.5��                          4                     5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                v       f?o     �                3.5��                          �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                          f?t     �               htype TRANSMISSOR is (DISPONIVEL, TRANSMITINDO, ESPERA); -- Declaração do tipo da máquina de ESTADOs     Bsignal ESTADO: TRANSMISSOR; -- Declaração da máquina de ESTADOs�               �signal PALAVRA_TRANSMITIR: std_logic_vector (9 downto 0) := "1111111111"; -- Vetor que guardará a palavra a ser enviada via serial     5��                          �                     �                          8                     �                          �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                          f?x     �               F    signal ESTADO: TRANSMISSOR; -- Declaração da máquina de ESTADOs5��                        �                    5�_�                       	    ����                                                                                                                                                                                                                                                                                                                                                          f?�     �               l    type TRANSMISSOR is (DISPONIVEL, TRANSMITINDO, ESPERA); -- Declaração do tipo da máquina de ESTADOs  5��       	              
   A             
       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                          f?�     �               k    type transmiter is (DISPONIVEL, TRANSMITINDO, ESPERA); -- Declaração do tipo da máquina de ESTADOs  5��              
       	   P      
       	       5�_�                       #    ����                                                                                                                                                                                                                                                                                                                                                          f?�     �               j    type transmiter is (available, TRANSMITINDO, ESPERA); -- Declaração do tipo da máquina de ESTADOs  5��       #                 [                    �       #                 [                    �       #                 [                    5�_�                       ,    ����                                                                                                                                                                                                                                                                                                                                                          f?�     �               e    type transmiter is (available, sending, ESPERA); -- Declaração do tipo da máquina de ESTADOs  5��       ,                 d                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                          f?�     �               �    signal PALAVRA_TRANSMITIR: std_logic_vector (9 downto 0) := "1111111111"; -- Vetor que guardará a palavra a ser enviada via serial     5��                        �                    �       !                  �                     �                          �                     �                        �                    �       !                  �                     �                          �                     �                     
   �             
       �              
       
   �      
       
       �              
          �      
              �                     
   �             
       5�_�                       )    ����                                                                                                                                                                                                                                                                                                                                                          f?�     �               �    signal PALAVRA_TRANSMITIR: bit_vector (9 downto 0) := "1111111111"; -- Vetor que guardará a palavra a ser enviada via serial     5��       )                  �                     5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                                          f?�     �               �    signal PALAVRA_TRANSMITIR: bit_vector(9 downto 0) := "1111111111"; -- Vetor que guardará a palavra a ser enviada via serial     5��       *                 �                    �       +                  �                     �       *                 �                    �       *                 �                    �       *                 �                    5�_�                       M    ����                                                                                                                                                                                                                                                                                                                                                          f?�     �               �    signal PALAVRA_TRANSMITIR: bit_vector(WIDTH-1 downto 0) := "1111111111"; -- Vetor que guardará a palavra a ser enviada via serial     5��       M       >           �      >               5�_�                       L    ����                                                                                                                                                                                                                                                                                                                                                          f?�     �               M    signal PALAVRA_TRANSMITIR: bit_vector(WIDTH-1 downto 0) := "1111111111"; 5��       L                  �                     5�_�                       2    ����                                                                                                                                                                                                                                                                                                                                                          f?�     �               c    type transmiter is (available, sending, idle); -- Declaração do tipo da máquina de ESTADOs  5��       2       1           *      1               5�_�                           ����                                                                                                                                                                                                                                                                                                                                                          f?�     �               E    signal state: TRANSMISSOR; -- Declaração da máquina de ESTADOs5��                        =                    �                         ?                     �                         >                     �                     
   =             
       �              
          =      
              �                     
   =             
       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                          f?�    �               L    signal PALAVRA_TRANSMITIR: bit_vector(WIDTH-1 downto 0) := "1111111111";5��                        �                    5�_�                       0    ����                                                                                                                                                                                                                                                                                                                                                          f�8     �               >    signal word: bit_vector(WIDTH-1 downto 0) := "1111111111";5��       0                  �                     �       /                  �                     �       -                  �                     5�_�                       ,    ����                                                                                                                                                                                                                                                                                                                                                          f�H     �                2    type transmiter is (available, sending, idle);5��                          �      3               5�_�                       ,    ����                                                                                                                                                                                                                                                                                                                                                          f�I     �             �             5��                          �              3       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                          f�K     �             5��                          �                     �                          �                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                                          f�.     �                   5��                         g                     5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                                          f�>     �                   OI5��                        h                    5�_�       "           !          ����                                                                                                                                                                                                                                                                                                                                                          f�f     �                   Oi5��                        g                    5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                                                          f�4     �                   OI5��                         g                     �                         f                     �                         e                     �                         d                     �                          c                     5�_�   "   $           #           ����                                                                                                                                                                                                                                                                                                                                                          f�W     �                5��                          c                     5�_�   #   &           $           ����                                                                                                                                                                                                                                                                                                                                                          f�_     �               i5��                         c                    �                         f                     �                         e                     �                         d                     �                          c                     5�_�   $   '   %       &          ����                                                                                                                                                                                                                                                                                                                                                          f�     �               2    type transmiter is (available, sending, idle);5��              	          �      	              5�_�   &   (           '      +    ����                                                                                                                                                                                                                                                                                                                                                          f�     �               1    type transmiter is (starting, sending, idle);5��       +                 �                    5�_�   '   )           (      -    ����                                                                                                                                                                                                                                                                                                                                                          f��     �                .    signal word: bit_vector(WIDTH-1 downto 0);5��                          �      /               5�_�   (   *           )      ;    ����                                                                                                                                                                                                                                                                                                                                                          f��     �             �             5��                          -              /       5�_�   )   +           *          ����                                                                                                                                                                                                                                                                                                                                                          f��     �                D    signal state: transmiter; -- Declaração da máquina de ESTADOs5��                          �      E               5�_�   *   ,           +           ����                                                                                                                                                                                                                                                                                                                                                          f��     �             �             5��                          �              E       5�_�   +   -           ,           ����                                                                                                                                                                                                                                                                                                                                         8       v   8    f�     �      -          �             5��                          l                     �                        p              �      5�_�   ,   .           -           ����                                                                                                                                                                                                                                                                                                                                       ,                   f�      �      -   .          if rising_edge(Clk) then           if nRst = '0' then   #            State <= <reset_state>;           else               case State is   $                when <state_name> =>   5                    <set_outputs_for_this_state_here>   <                    if <state_change_condition_is_true> then   3                        State <= <next_state_name>;                       end if;                   ...               end case;           end if;       end if;   end process;�         .      begin5��                          �                     �                          �                     �                          �                     �                          �                     �                           �                     �    !                                           �    "                      !                     �    #                      J                     �    $                      �                     �    %                      �                     �    &                      �                     �    '                                           �    (                      5                     �    )                      O                     �    *                      c                     �    +                      s                     5�_�   -   /           .          ����                                                                                                                                                                                                                                                                                                                                       ,                   f�'     �         .          process(Clk) is5��                        x                    �                        x                    �                        x                    �                        x                    5�_�   .   0           /          ����                                                                                                                                                                                                                                                                                                                                                V       f�-     �         .               if rising_edge(Clk) then5��                        �                    �                        �                    �                        �                    �                        �                    5�_�   /   1           0          ����                                                                                                                                                                                                                                                                                                                                                V       f�1     �          .                  if nRst = '0' then5��                        �                    �                        �                    �                        �                    �                        �                    �                        �                    5�_�   0   2           1           ����                                                                                                                                                                                                                                                                                                                                                V       f�:     �      !   .      '                State <= <reset_state>;5��                        �                    5�_�   1   3           2           ����                                                                                                                                                                                                                                                                                                                                                V       f�F     �      !   .      '                state <= <reset_state>;5��                        �                    5�_�   2   5           3           ����                                                                                                                                                                                                                                                                                                                                                V       f�J     �      !   .                      state <= idle;5��                         �                     5�_�   3   6   4       5   "       ����                                                                                                                                                                                                                                                                                                                                                V       f�R     �   !   #   .                      case State is5��    !                                        �    !                     "                     �    !                     !                     �    !                                           �    !                                        �    !                                        �    !                                        5�_�   5   7           6   '        ����                                                                                                                                                                                                                                                                                                                            #          '          V       f��     �   '   -   .    �   '   (   .    5��    '                      $              �       5�_�   6   8           7   ,       ����                                                                                                                                                                                                                                                                                                                            #          '          V       f��     �   ,   2   3    �   ,   -   3    5��    ,                                     �       5�_�   7   9           8   2       ����                                                                                                                                                                                                                                                                                                                            #          '          V       f��     �   1   2                              ...5��    1                                           5�_�   8   :           9   #       ����                                                                                                                                                                                                                                                                                                                            #          '          V       f��     �   "   $   7      (                    when <state_name> =>5��    "                    A                    5�_�   9   ;           :   $       ����                                                                                                                                                                                                                                                                                                                            #          '          V       f��     �   #   %   7      9                        <set_outputs_for_this_state_here>5��    #          !          a      !              �    #                     d                     �    #                     c                     �    #                     b                     �    #                    a                    �    #                    a                    �    #                    a                    5�_�   :   <           ;   $   #    ����                                                                                                                                                                                                                                                                                                                            #          '          V       f�      �   #   %   7      #                        tx_done <= 5��    #   #                  l                     5�_�   ;   =           <   $   $    ����                                                                                                                                                                                                                                                                                                                            #          '          V       f�      �   #   %   7      %                        tx_done <= ''5��    #   $                  m                     5�_�   <   >           =   $   &    ����                                                                                                                                                                                                                                                                                                                            #          '          V       f�     �   #   %   7      &                        tx_done <= '1'5��    #   &                  o                     5�_�   =   ?           >   $   &    ����                                                                                                                                                                                                                                                                                                                            #          '          V       f�     �   $   &   8                              �   $   &   7    5��    $                      q                     �    $                     �                     �    $                     �                     �    $                     �                     �    $                 
   �             
       �    $          
          �      
              �    $                 
   �             
       �    $   !                  �                     �    $                      �                     �    $                    �                    5�_�   >   @           ?   %   $    ����                                                                                                                                                                                                                                                                                                                            #          (          V       f�     �   $   &   8      $                        serial_o <= 5��    $   $                  �                     5�_�   ?   A           @   %   %    ����                                                                                                                                                                                                                                                                                                                            #          (          V       f�     �   $   &   8      &                        serial_o <= ''5��    $   %                  �                     5�_�   @   B           A   %   '    ����                                                                                                                                                                                                                                                                                                                            #          (          V       f�     �   $   &   8      '                        serial_o <= '1'5��    $   '                  �                     5�_�   A   C           B   &       ����                                                                                                                                                                                                                                                                                                                            #          (          V       f�     �   %   '   8      @                        if <state_change_condition_is_true> then5��    %                     �                     �    %                     �                     �    %                    �                    �    %                     �                     �    %                     �                     �    %                    �                    �    %                    �                    �    %                    �                    5�_�   B   D           C          ����                                                                                                                                                                                                                                                                                                                               -                 v   I    f�H     �         9          �         8    5��                          \                     �                         `                     �                         k                     �                        j                    �                        q                    5�_�   C   E           D   '   #    ����                                                                                                                                                                                                                                                                                                                               -                 v   I    f�b     �   &   (   9      (                        if state =  then5��    &   #                  �                     �    &   &                  �                     �    &   %                  �                     �    &   $                  �                     �    &   #                 �                    �    &   #                 �                    �    &   #              
   �             
       �    &   ,                 �                    �    &   ,                  �                     5�_�   D   F           E   '       ����                                                                                                                                                                                                                                                                                                                               -                 v   I    f�i     �   &   (   9      1                        if state = stopping  then5��    &                     �                     5�_�   E   G           F   '       ����                                                                                                                                                                                                                                                                                                                               -                 v   I    f�k     �   &   (   9      2                        if (state = stopping  then5��    &                     �      3       4       5�_�   F   H           G   '   -    ����                                                                                                                                                                                                                                                                                                                               -                 v   I    f�m     �   &   (   9      3                        if (state = stopping)  then5��    &   -                  �                     5�_�   G   I           H   '   2    ����                                                                                                                                                                                                                                                                                                                               -                 v   I    f�p     �   &   (   9      8                        if (state = stopping) and   then5��    &   2                  �                     5�_�   H   J           I   '   2    ����                                                                                                                                                                                                                                                                                                                               -                 v   I    f�s     �   &   (   9      7                        if (state = stopping) and  then5��    &   2                  �                     �    &   5                  �                     �    &   4                  �                     �    &   3                  �                     �    &   2                 �                    �    &   2                 �                    �    &   2                 �                    5�_�   I   K           J   '   =    ����                                                                                                                                                                                                                                                                                                                               -                 v   I    f�v     �   &   (   9      B                        if (state = stopping) and finished =  then5��    &   =                  �                     5�_�   J   L           K   '   >    ����                                                                                                                                                                                                                                                                                                                               -                 v   I    f�w     �   &   (   9      D                        if (state = stopping) and finished = '' then5��    &   >                  �                     5�_�   K   M           L   (   %    ����                                                                                                                                                                                                                                                                                                                               -                 v   I    f��     �   '   )   9      7                            State <= <next_state_name>;5��    '   %                                     �    '   &                                        �    '   %                                     �    '   %                                     �    '   %                                     5�_�   L   N           M   '       ����                                                                                                                                                                                                                                                                                                                            '          '   1       v   1    f��     �   &   (   9      E                        if (state = stopping) and finished = '1' then5��    &                     �                     5�_�   M   O           N   '       ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f��     �   &   (   9      .                        if finished = '1' then5��    &                    �                    �    &                     �                     �    &                    �                    �    &   !                  �                     �    &                      �                     �    &                     �                     �    &                     �                     �    &                     �                     �    &                     �                     �    &                    �                    �    &                     �                     �    &                     �                     �    &                     �                     �    &                     �                     �    &                    �                    �    &                    �                    �    &                    �                    5�_�   N   P           O   '   #    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f��     �   &   (   9      (                        if tx_go =  then5��    &   #                  �                     5�_�   O   Q           P   '   $    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f��     �   &   (   9      *                        if tx_go = '' then5��    &   $                  �                     5�_�   P   R           Q   (       ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f��     �   '   )   9      *                            State <= idle;5��    '                    �                    5�_�   Q   S           R           ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�     �      !   9                  if reset = '0' then5��                        �                    5�_�   R   T           S   *       ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�     �   )   +   9      (                    when <state_name> =>5��    )                    D                    �    )                     G                     �    )                     F                     �    )                     E                     �    )                    D                    �    )                    D                    �    )                    D                    5�_�   S   U           T   +       ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�(     �   *   ,   9      9                        <set_outputs_for_this_state_here>5��    *          !          h      !              �    *                     i                     �    *                    h                    �    *                     l                     �    *                     k                     �    *                     j                     �    *                     i                     �    *                    h                    �    *                     n                     �    *                     m                     �    *                     l                     �    *                     k                     �    *                     j                     �    *                     i                     �    *                    h                    �    *                    h                    �    *                    h                    5�_�   T   V           U   +   #    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�0     �   *   ,   9      #                        tx_done <= 5��    *   #                  s                     5�_�   U   W           V   +   $    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�0     �   *   ,   9      %                        tx_done <= ''5��    *   $                  t                     5�_�   V   X           W   +   &    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�2     �   +   -   :                               serial_o�   *   -   9      &                        tx_done <= '0'5��    *   &                  v                     �    *   '                 w                     �    +                     �                     �    +                     �                     �    +                     �                     �    +                     �                     �    +                    �                    �    +                     �                     �    +                     �                     �    +                     �                     �    +                     �                     �    +                     �                     �    +                     �                     �    +                     �                     �    +                    �                    �    +                    �                    �    +                    �                    5�_�   W   Y           X   ,   #    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�9     �   +   -   :      #                        serial_o <=5��    +   #                  �                     5�_�   X   Z           Y   ,   $    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�:     �   +   -   :      $                        serial_o <= 5��    +   $                  �                     5�_�   Y   [           Z   ,   %    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�:     �   +   -   :      &                        serial_o <= ''5��    +   %                  �                     5�_�   Z   \           [   ,   '    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�;     �   +   -   :      '                        serial_o <= '0'5��    +   '                  �                     5�_�   [   ]           \   -       ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�?     �   ,   .   :      @                        if <state_change_condition_is_true> then5��    ,                      �                      5�_�   \   ^           ]   -       ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�F     �   ,   -                                   if  then5��    ,                      �      !               5�_�   ]   _           ^   .       ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�G     �   -   .                                  end if;5��    -                      �                      5�_�   ^   `           _   -       ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�H     �   ,   .   8      7                            State <= <next_state_name>;5��    ,                     �                     �    ,                     �                     �    ,                     �                     �    ,                     �                     5�_�   _   a           `   -       ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�L     �   ,   .   8      3                        State <= <next_state_name>;5��    ,                    �                    5�_�   `   b           a   -   !    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�P     �   ,   .   8      3                        state <= <next_state_name>;5��    ,   !                 �                    �    ,   #                  �                     �    ,   "                  �                     �    ,   !                 �                    �    ,   #                  �                     �    ,   "                  �                     �    ,   !                 �                    �    ,   !                 �                    �    ,   !                 �                    5�_�   a   c           b   -   '    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�Y     �   ,   .   9                              �   ,   .   8    5��    ,                      �                     �    ,                     �                     �    ,                     �                     �    ,                     �                     �    ,                     �                     �    ,                    �                    �    ,                    �                    �    ,                    �                    5�_�   b   d           c   -   $    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�_     �   ,   .   9      $                        finished <= 5��    ,   $                  �                     5�_�   c   e           d   -   %    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�`     �   ,   .   9      &                        finished <= ''5��    ,   %                  �                     5�_�   d   f           e   -   '    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�a     �   ,   .   9      '                        finished <= '0'5��    ,   '                  �                     5�_�   e   g           f   (   %    ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�x     �   '   )   9      *                            state <= idle;5��    '   %                                     �    '   '                                       �    '   &                                       �    '   %                                     �    '   %                                     �    '   %                                     5�_�   f   h           g   /       ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f��     �   .   0   9      (                    when <state_name> =>5��    .                                        �    .                                          �    .                                          �    .                                        �    .                                        �    .                                        5�_�   g   i           h          ����                                                                                                                                                                                                                                                                                                                            '          '   (       v   (    f�F     �         :          �         9    5��                          v                     �                         z                     �                         �                     �                        �                    5�_�   h   j           i          ����                                                                                                                                                                                                                                                                                                                            (          (   (       v   (    f�[     �         :          signal stopped_bits:5��                      	   �              	       5�_�   i   k           j   .        ����                                                                                                                                                                                                                                                                                                                            (          (   (       v   (    f�|     �   -   .          (                        finished <= '0';5��    -                      �      )               5�_�   j   l           k   .        ����                                                                                                                                                                                                                                                                                                                            (          (   (       v   (    f�~     �   -   /   9    �   .   /   9    5��    -                      �              )       5�_�   k   m           l   .       ����                                                                                                                                                                                                                                                                                                                            (          (   (       v   (    f�     �   -   /   :      (                        finished <= '0';5��    -                    �                    �    -                     �                     �    -                     �                     �    -                     �                     �    -                    �                    �    -                     �                     �    -                     �                     �    -                     �                     �    -                     �                     �    -                     �                     �    -                     �                     �    -                     �                     �    -                    �                    �    -   #                  �                     �    -   "                  �                     �    -   !                  �                     �    -                      �                     �    -                     �                     �    -                     �                     �    -                     �                     �    -                     �                     �    -                     �                     �    -                     �                     �    -                     �                     �    -                    �                    �    -                    �                    �    -                    �                    5�_�   l   n           m   .   '    ����                                                                                                                                                                                                                                                                                                                            (          (   (       v   (    f��     �   -   /   :      ,                        stopped_bits <= '0';5��    -   '                 �                    �    -   '                 �                    5�_�   m   o           n   .   (    ����                                                                                                                                                                                                                                                                                                                            (          (   (       v   (    f��     �   -   .          *                        stopped_bits <= 0;5��    -                      �      +               5�_�   n   p           o   '   '    ����                                                                                                                                                                                                                                                                                                                            (          (   (       v   (    f��    �   '   )   9    �   '   (   9    5��    '                      �              +       5�_�   o   q           p      =    ����                                                                                                                                                                                                                                                                                                                                                             f�     �         :      D    signal state: transmiter; -- Declaração da máquina de ESTADOs5��       =                 $                    5�_�   p   r           q   4        ����                                                                                                                                                                                                                                                                                                                            0   "       4          V   @    f��     �   4   :   :    �   4   5   :    5��    4                                    �       5�_�   q   s           r          ����                                                                                                                                                                                                                                                                                                                            0   "       4          V   @    f��     �         @          �         ?    5��                          v                     �                         z                     �                         �                     �                        �                    5�_�   r   t           s          ����                                                                                                                                                                                                                                                                                                                            1   "       5          V   @    f��     �         @          signal bits_sent: nat5��                         �                     5�_�   s   u           t          ����                                                                                                                                                                                                                                                                                                                            1   "       5          V   @    f��     �         @          signal bits_sent: nat[]5��                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    5�_�   t   v           u   )       ����                                                                                                                                                                                                                                                                                                                            1   "       5          V   @    f��     �   )   +   @    �   )   *   @    5��    )                                     +       5�_�   u   w           v   *       ����                                                                                                                                                                                                                                                                                                                            2   "       6          V   @    f��     �   )   +   A      *                        stopped_bits <= 0;5��    )                    8                    �    )                    8                    �    )                 	   8             	       �    )          	       	   8      	       	       �    )          	          8      	              �    )                 	   8             	       5�_�   v   x           w          ����                                                                                                                                                                                                                                                                                                                            2   "       6          V   @    f�q     �          A    5��                                                  5�_�   w   y           x           ����                                                                                                                                                                                                                                                                                                                            3   "       7          V   @    f�r    �       '   B    �         B    5��                    &                       �      5�_�   x   z           y   :       ����                                                                                                                                                                                                                                                                                                                            Y   "       ]          V   @    f��     �   <   >   k          end component�   ;   >   j          component counter_generic�   :   =   i          �   :   <   h    5��    :                      8                     �    :                      8                     �    :                      8                     �    :                     8                     �    ;                     =                     �    ;                     K                     �    ;                     J                     �    ;                     I                     �    ;                     H                     �    ;                    G                    �    ;                    G                    �    ;                    G                    �    ;                     X                     �    ;                     W                     �    ;                     V                     �    ;                    V                     �    <                     W                    �    <   
                  a                     �    <   	                  `                     �    <                    _                    �    <                     W                    �    <                     _                     �    <   
                  a                     �    <   	                  `                     �    <                 	   _             	       �    <          	          _      	              �    <                 
   _             
       �    <                    h                    5�_�   y   {           z   <        ����                                                                                                                                                                                                                                                                                                                                                V       f��     �   <   E   k    �   <   =   k    5��    <                      W              �       5�_�   z   |           {   =       ����                                                                                                                                                                                                                                                                                                                            =          D                 f��     �   =   E   s              MAX_COUNT: natural       );   
    port (   J        clk, rst, start: in bit;                            -- Clock input           done: out bit;   B        count : out natural       -- 6-bit count output (64 steps)       );�   <   >   s          generic(5��    <                     [                     �    =                     l                     �    >                     �                     �    ?                     �                     �    @                     �                     �    A                     �                     �    B                                          �    C                     V                     5�_�   {   }           |   O       ����                                                                                                                                                                                                                                                                                                                            =          D                 f�     �   Q   S   v              generic�   P   S   u      !    count_signal: counter_generic�   O   R   t          �   O   Q   s    5��    O                      �                     �    O                      �                     �    O                      �                     �    O                     �                     �    P                  	   �              	       �    P                     �                     �    P                     �                     �    P   
                 �                    �    P                     �                     �    P                     �                     �    P   
                 �                    �    P                     �                     �    P   
                 �                    �    P                     �                     �    P                     �                     �    P                     �                     �    P                     �                     �    P                    �                    �    P                    �                    �    P                    �                    �    P   !                  �                     �    P   !                 �                     �    Q                     �                     �    Q                    �                    �    Q                    �                    �    Q                    �                    5�_�   |   ~           }   R       ����                                                                                                                                                                                                                                                                                                                            =          D                 f�     �   Q   S   v              generic map5��    Q                     �                     5�_�   }              ~   R       ����                                                                                                                                                                                                                                                                                                                            =          D                 f�      �   Q   S   v              generic map()5��    Q                     �                     �    Q                    �                    �    Q                    �                    �    Q                    �                    �    Q                     �                     �    Q                     �                     5�_�   ~   �              R       ����                                                                                                                                                                                                                                                                                                                            =          D                 f�'     �   R   T   w              port�   Q   T   v              generic map(WIDTH)5��    Q                    �              	       �    R                     �                     �    R                    �                    �    R                    �                    �    R                    �                    5�_�      �           �   S       ����                                                                                                                                                                                                                                                                                                                            =          D                 f�*     �   R   T   w              port map5��    R                     �                     5�_�   �   �           �   S       ����                                                                                                                                                                                                                                                                                                                            =          D                 f�/     �   R   T   w              port map()5��    R                     �                     �    R                    �                    �    R                    �                    �    R                 
   �             
       �    R                    �                    �    R                    �                    �    R                 	   �             	       5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            =          D                 f�@     �   K   L              signal bits_sent: natural;5��    K                      <                     5�_�   �   �           �   L        ����                                                                                                                                                                                                                                                                                                                            =          D                 f�A     �   K   L          !    signal stopped_bits: natural;5��    K                      <      "               5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                            =          D                 f�D     �   J   L   u          signal finished: bit;5��    J                     5                     5�_�   �   �           �   Q   !    ����                                                                                                                                                                                                                                                                                                                            =          D                 f�a     �   P   R   u      "        port map(clock, reset, , )5��    P   !                  �                     �    P   !                 �                    �    P   !                 �                    �    P   !                 �                    �    P   2                 �                    �    P   =                 �                    5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                            =          D                 f��     �   K   M   v          �   K   M   u    5��    K                      C                     �    K                     G                     5�_�   �   �           �   L   
    ����                                                                                                                                                                                                                                                                                                                            =          D                 f��     �   K   M   v          signal �   L   M   v    5��    K                     N                     5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            =          D                 f��     �   K   M   v          signal signal_bits_sent5��    K                     ^                     �    K                      c                     �    K                     b                     �    K                     a                     �    K                    `                    �    K                    `                    �    K                    `                    5�_�   �   �           �   L   $    ����                                                                                                                                                                                                                                                                                                                            =          D                 f��     �   K   M   v      $    signal signal_bits_sent: natural5��    K   $                  g                     5�_�   �   �   �       �   K       ����                                                                                                                                                                                                                                                                                                                            =          D                 f��     �   J   L   v    5��    J                      "                     5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                            =          D                 f��     �   J   L   w          5��    J                     &                     5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                            =          D                 f��     �   J   M   w          []5��    J                     &                     �    J                     &                     �    J                    &                     �    K                     +                     5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            =          D                 f��     �   S   U   x      C        port map(clock, reset, , finished_signal, signal_bits_sent)5��    S                     �                     �    S                    �                    �    S                    �                    �    S                    �                    5�_�   �   �           �   T   N    ����                                                                                                                                                                                                                                                                                                                            =          D                 f��     �   S   U   x      N        port map(clock, reset, send_signal, finished_signal, signal_bits_sent)5��    S   N                  "                     5�_�   �   �           �   T        ����                                                                                                                                                                                                                                                                                                                            R           T   N       V   N    f�     �   T   V   x    5��    T                      $              	       �    T                      $                     5�_�   �   �           �   U        ����                                                                                                                                                                                                                                                                                                                            R           T   N       V   N    f�     �   U   Y   y    �   U   V   y    5��    U                      %              �       5�_�   �   �           �   V   
    ����                                                                                                                                                                                                                                                                                                                            R           T   N       V   N    f�     �   U   W   |      !    count_signal: counter_generic5��    U   
                 /                    �    U                     3                     5�_�   �   �           �   W       ����                                                                                                                                                                                                                                                                                                                            R           T   N       V   N    f�     �   V   X   |              generic map(WIDTH)5��    V                    Y                    �    V                 	   Y             	       �    V          	          Y      	              �    V                 	   Y             	       5�_�   �   �           �   N        ����                                                                                                                                                                                                                                                                                                                            L          N          V       f�!     �   N   P   |    5��    N                      �                     �    N                      �                     5�_�   �   �           �   O        ����                                                                                                                                                                                                                                                                                                                            L          N          V       f�!     �   O   S   }    �   O   P   }    5��    O                      �              d       5�_�   �   �           �   P       ����                                                                                                                                                                                                                                                                                                                            L          N          V       f�(     �   O   Q   �          signal send_signal: bit;5��    O                    �                    5�_�   �   �           �   Q       ����                                                                                                                                                                                                                                                                                                                            L          N          V       f�+     �   P   R   �           signal finished_signal: bit;5��    P                    �                    5�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                            R          R          v       f�1     �   Q   S   �      %    signal signal_bits_sent: natural;5��    Q                    �                    5�_�   �   �           �   \        ����                                                                                                                                                                                                                                                                                                                            \          \          V       f�>     �   [   ]   �      O        port map(clock, reset, send_signal, finished_signal, signal_bits_sent);5��    [   $                 �                    �    [   3                 �                    �    [   9                 �                    5�_�   �   �           �   L        ����                                                                                                                                                                                                                                                                                                                            L          \          V       f�,     �   [   ]          I        port map(clock, reset, send_stop, finished_stop, stop_bits_sent);�   W   Y          O        port map(clock, reset, send_signal, finished_signal, signal_bits_sent);�   O   Q              signal send_stop: bit;�   K   M   �          signal send_signal: bit;5��    K                    2                    �    O                    �                    �    W                    T                    �    [                    �                    5�_�   �   �   �       �   M        ����                                                                                                                                                                                                                                                                                                                            \           M           V        f�Y    �   [   ]          J        port map(clock, reset, start_stop, finished_stop, stop_bits_sent);�   W   Y          P        port map(clock, reset, start_signal, finished_signal, signal_bits_sent);�   P   R              signal finished_stop: bit;�   L   N   �           signal finished_signal: bit;5��    L                    P                    �    P                    �                    �    W   -                 Z                    �    [   +                 �                    5�_�   �   �           �   f        ����                                                                                                                                                                                                                                                                                                                                                             f��     �   e   g   �    5��    e                      �	                     �    e                      �	                     5�_�   �   �           �   f        ����                                                                                                                                                                                                                                                                                                                                                             f��     �   e   f           5��    e                      �	                     5�_�   �   �           �   g       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   g   j   �                              �   g   i   �    5��    g                      4
                     �    g                      4
                     �    g                     4
                     �    h                  
   M
              
       5�_�   �   �           �   l   !    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   k   m   �    5��    k                      �
                     �    k                      �
                     5�_�   �   �           �   j       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   i   k   �      *                        stopped_bits <= 0;5��    i                    p
                    �    i                    r
                    �    i                    p
                    �    i                    p
                    �    i                 
   p
             
       �    i          
          p
      
              �    i                    p
                    �    i                    p
                    �    i                    p
                    5�_�   �   �           �   j   )    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   i   k   �      *                        start_signal <= 0;5��    i   (                  �
                     5�_�   �   �           �   j   (    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   i   k   �      )                        start_signal <= ;5��    i   (                  �
                     5�_�   �   �           �   j   )    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   i   k   �      +                        start_signal <= '';5��    i   )                  �
                     5�_�   �   �           �   j   )    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   j   l   �    �   j   k   �    5��    j                      �
              -       5�_�   �   �           �   l       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   k   l          '                        bits_sent <= 0;5��    k                      �
      (               5�_�   �   �           �   k       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   j   l   �      ,                        start_signal <= '1';5��    j                    �
                    5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   K   M   �          signal start_signal: bit;5��    K                     2                     5�_�   �   �           �   P   
    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   O   Q   �          signal start_stop: bit;�   P   Q   �    5��    O                     �                     5�_�   �   �           �   P       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   O   Q   �      '    signal start_signalstart_stop: bit;5��    O                     �                     5�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   L   N   �          signal done_signal: bit;5��    L                     D                     5�_�   �   �           �   Q   
    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   P   R   �          signal done_stop: bit;�   Q   R   �    5��    P                     �                     5�_�   �   �           �   Q       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   P   R   �      %    signal done_signaldone_stop: bit;5��    P                     �                     5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   M   O   �      %    signal signal_bits_sent: natural;5��    M                     V                     5�_�   �   �           �   R   
    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   Q   S   �      #    signal stop_bits_sent: natural;�   R   S   �    5��    Q                     �                     5�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   Q   S   �      3    signal signal_bits_sentstop_bits_sent: natural;5��    Q                     �                     5�_�   �   �           �   L        ����                                                                                                                                                                                                                                                                                                                                                             f�      �   K   L              signal : bit;       signal : bit;       signal : natural;    5��    K                      '      ;               5�_�   �   �           �   L   (    ����                                                                                                                                                                                                                                                                                                                                                             f�     �   K   M         )    signal start_signal, start_stop: bit;5��    K   (                  O                     5�_�   �   �           �   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             f�     �   K   M         -    signal start_signal, start_stop: bit := ;5��    K   ,                  S                     5�_�   �   �           �   L   -    ����                                                                                                                                                                                                                                                                                                                                                             f�     �   K   M         /    signal start_signal, start_stop: bit := '';5��    K   -                  T                     5�_�   �   �           �   H       ����                                                                                                                                                                                                                                                                                                                                                             f�     �   G   I         D    signal state: transmiter; -- Declaração da máquina de estados5��    G                     �                     �    G                     �                     �    G                    �                    5�_�   �   �           �   L   (    ����                                                                                                                                                                                                                                                                                                                                                             f�     �   K   M         0    signal start_signal, start_stop: bit := '0';5��    K   (                  W                     5�_�   �   �           �   f   )    ����                                                                                                                                                                                                                                                                                                                                                             f�,     �   e   g         ,                        start_signal <= '1';5��    e   )                 T
                    5�_�   �   �           �   g   '    ����                                                                                                                                                                                                                                                                                                                                                             f�-     �   f   h         *                        start_stop <= '1';5��    f   '                 
                    5�_�   �   �   �       �   n   !    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�a     �   n   p       5��    n                      u                     �    n                      u                     5�_�   �   �           �   o        ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�a     �   o   s   �    �   o   p   �    5��    o                      v              {       5�_�   �   �           �   s       ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�d     �   r   t   �    5��    r                      �                     �    r                      �                     5�_�   �   �           �   q   )    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�i     �   p   r   �      ,                        start_signal <= '0';5��    p   )                 �                    5�_�   �   �           �   r   '    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�j     �   q   s   �      *                        start_stop <= '0';5��    q   '                 �                    5�_�   �   �   �       �   r   '    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f��     �   r   t   �                              �   r   t   �    5��    r                      �                     �    r                     	                     �    r                     
                     �    r                    	                    �    r                    	                    �    r                    	                    5�_�   �   �           �   g       ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f��     �   g   i   �                              �   g   i   �    5��    g                      �
                     �    g                     �
                     �    g                     �
                     �    g                    �
                    �    g                    �
                    �    g                 
   �
             
       �    g   !                  �
                     �    g                     �
                    �    g                     �
                    �    g                     �
                    �    g                     �
                    5�_�   �   �           �   h        ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f��     �   g   i   �      -                        word <= others => '0'5��    g                      �
                     5�_�   �   �           �   h   !    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f��     �   g   i   �      .                        word <= (others => '0'5��    g                     �
      /       0       5�_�   �   �           �   h   -    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f��     �   g   i   �      /                        word <= (others => '0)'5��    g   -                  �
                     5�_�   �   �           �   h   -    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f��     �   g   i   �      .                        word <= (others => '0'�   h   i   �    5��    g   .                  �
                     5�_�   �   �           �   h   /    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f��     �   g   i   �      /                        word <= (others => '0')5��    g   /                  �
                     5�_�   �   �           �   t       ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f��     �   s   u   �                              word <=5��    s                     A                     �    s   !                  C                     �    s                      B                     5�_�   �   �           �   t        ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f��     �   s   u   �                               word <= 5��    s                      B                     5�_�   �   �           �   z       ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�#     �   y   {   �      7                            State <= <next_state_name>;5��    y                    .                    5�_�   �   �           �   z   %    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�,     �   y   {   �      7                            state <= <next_state_name>;5��    y   %                 7                    5�_�   �   �           �   y       ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�2     �   x   z   �      @                        if <state_change_condition_is_true> then5��    x                      �                      5�_�   �   �           �   y       ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�O     �   x   z   �                               if  then5��    x                     �                     �    x                    �                    �    x                 	   �             	       �    x          	          �      	              �    x                    �                    �    x                    �                    �    x                    �                    5�_�   �   �           �   y   *    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�a     �   x   z   �      /                        if done_signal /=  then5��    x   *                  �                     5�_�   �   �           �   y   +    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�b     �   x   z   �      1                        if done_signal /= '' then5��    x   +                  �                     5�_�   �   �           �   x       ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�y     �   w   y   �      9                        <set_outputs_for_this_state_here>5��    w          !          �      !              �    w                     �                     �    w                     �                     �    w                    �                    �    w                    �                    �    w                    �                    5�_�   �   �           �   x   "    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f��     �   x   z   �    5��    x                      �                     �    x                     �                    �    x                      �                     5�_�   �   �           �   x   #    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f��     �   w   y   �      #                        serial_o <=5��    w   #                  �                     �    w   %                  �                     �    w   $                 �                    �    w   $                 �                    �    w   $                 �                    �    w   (                  �                     5�_�   �   �           �   x   (    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�X     �   w   y   �      (                        serial_o <= word5��    w   (                  �                     5�_�   �   �           �   x   )    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�Z     �   w   y   �      *                        serial_o <= word()5��    w   )                  �                     �    w   )                 �                    �    w   )                 �                    �    w   )                 �                    �    w   1                 �                    �    w   1                  �                     5�_�   �   �           �   x   0    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�u     �   w   y   �      2                        serial_o <= word(WIDTH-1-)�   x   y   �    5��    w   1                  �                     5�_�   �   �           �   x   B    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f�w     �   w   y   �      B                        serial_o <= word(WIDTH-1-signal_bits_sent)5��    w   B                  �                     5�_�   �   �           �   |        ����                                                                                                                                                                                                                                                                                                                f   '       z   1       |          V   B    f     �   |   �   �    �   |   }   �    5��    |                      ]              �       5�_�   �   �           �   z   '    ����                                                                                                                                                                                                                                                                                                                f   '       z   1       |          V   B    f     �   y   {   �      2                        if done_signal /= '1' then5��    y   '                                       5�_�   �   �           �   }   '    ����                                                                                                                                                                                                                                                                                                                f   '       z   1       |          V   B    f     �   |   ~   �      2                        if done_signal /= '1' then5��    |   '                  �                     5�_�   �   �           �   }   *    ����                                                                                                                                                                                                                                                                                                                f   '       z   1       |          V   B    f     �   |   ~   �      1                        if done_signal = '1' then5��    |   *                 �                    5�_�   �   �           �   z   *    ����                                                                                                                                                                                                                                                                                                                f   '       z   1       |          V   B    f     �   y   {   �      1                        if done_signal = '1' then5��    y   *                                     5�_�   �   �           �   }   *    ����                                                                                                                                                                                                                                                                                                                f   '       z   1       |          V   B    f      �   |   ~   �      1                        if done_signal = '0' then5��    |   *                 �                    5�_�   �   �           �   ~   %    ����                                                                                                                                                                                                                                                                                                                f   '       z   1       |          V   B    f£     �   }      �      -                            state <= sending;5��    }   %                 �                    �    }   '                 �                    �    }   '                 �                    �    }   %                 �                    �    }   %                 �                    �    }   %                 �                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                f   '       z   1       |          V   B    f´     �      �   �      #                    when sending =>5��                        �                    �                        �                    �                        �                    �                        �                    5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                f   '       z   1       |          V   B    f¹     �   �   �   �    5��    �                      <                     �    �                      <                     5�_�   �   �   �       �   W       ����                                                                                                                                                                                                                                                                                                                f   '       z   1       |          V   B    f��     �   V   X   �              generic map(STOP_BITS)5��    V                     �                     5�_�   �   �           �   W        ����                                                                                                                                                                                                                                                                                                                f   '       z   1       |          V   B    f��     �   V   X   �               generic map(STOP_BITS+1)5��    V                   
   �              
       �    V   (                 �                    �    V   )                 �                    �    V   .              
   �             
       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                f   '       z   1       |          V   B    f�r     �   �   �   �      9                        <set_outputs_for_this_state_here>5��    �          !          4      !              5�_�   �   �           �   s       ����                                                                                                                                                                                                                                                                                                                f   '       z   1       |          V   B    fÛ     �   r   s          *                        start_stop <= '1';5��    r                            +               5�_�   �   �           �   }       ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    fé     �   }      �    �   }   ~   �    5��    }                      �              +       5�_�   �   �           �   ~       ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    fê     �   }      �      *                        start_stop <= '1';5��    }                     �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    fö     �   �   �   �                              if 5��    �                     ;                     �    �                     >                     �    �                     =                     �    �                     <                     �    �                    ;                    �    �   (                  H                     �    �   '                  G                     �    �   &                  F                     �    �   %                  E                     �    �   $                  D                     �    �   #                  C                     �    �   "                  B                     �    �   !                  A                     �    �                      @                     �    �                     ?                     �    �                     >                     �    �                     =                     �    �                     <                     �    �                    ;                    �    �                    ;                    �    �                    ;                    5�_�   �   �           �   �   -    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f��     �   �   �   �      $                            serial_o�   �   �   �      -                        if stop_bits_sent = 05��    �   -                  M                     �    �   2                  R                     �    �   2                 R                     �    �                     S                    �    �                     q                     �    �                     p                     �    �                    o                    �    �                    o                    �    �                    o                    5�_�   �   �           �   �   +    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f��     �   �   �   �      +                            serial_o <= bit5��    �   +                  ~                     5�_�   �   �           �   �   ,    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f��     �   �   �   �      -                            serial_o <= bit()5��    �   ,                                       5�_�   �   �           �   �   4    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�      �   �   �   �      5                            serial_o <= bit(unsigned)5��    �   4                  �                     5�_�   �   �           �   �   5    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�     �   �   �   �      7                            serial_o <= bit(unsigned())5��    �   5                  �                     �    �   5                 �                    �    �   5                 �                    �    �   5                 �                    5�_�   �   �           �   �   =    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�     �   �   �   �      =                            serial_o <= bit(unsigned(PARITY))5��    �   =                  �                     5�_�   �   �           �   �   >    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�%     �   �   �   �      $                            serial_o�   �   �   �      >                            serial_o <= bit(unsigned(PARITY));5��    �   >                 �                     �    �                     �                     �    �                     �                    �    �                     �                     �    �                     �                     �    �                    �                     �    �                     �                    �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    �    �   (                  �                     5�_�   �   �           �   �   (    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�-     �   �   �   �      (                            serial_o <= 5��    �   (                  �                     5�_�   �   �           �   �   )    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�-     �   �   �   �      *                            serial_o <= ''5��    �   )                  �                     5�_�   �   �           �   �   +    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�.     �   �   �   �      +                            serial_o <= '1'5��    �   +                  �                     �    �   ,                 �                     �    �                     �                     �    �                     �                    �    �                     �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�5     �   �   �   �                              �   �   �   �    5��    �                                            �    �                     8                     �    �                    ;                    �    �                    ;                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�K     �   �   �   �      @                        if <state_change_condition_is_true> then5��    �                     8                     �    �                    8                    �    �                    8                    �    �                 	   8             	       �    �          	       	   8      	       	       �    �          	          8      	              �    �                    8                    5�_�   �   �           �   |       ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�^     �   {   }   �      1                        if done_signal = '1' then5��    {           1           K      1               5�_�   �   �           �   |        ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�`     �   {   |           5��    {                      K                     5�_�   �   �           �   {       ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�b     �   z   |   �                              end if;5��    z                     C                     �    z                      +                     �    z                     +                    5�_�   �   �           �   �   '    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�i     �   �   �   �      +                        if done_stop = then5��    �   '                                       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�n     �   �   �   �      7                            State <= <next_state_name>;5��    �                    4                    5�_�   �   �           �   �   %    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�p     �   �   �   �      7                            state <= <next_state_name>;5��    �   %                 =                    �    �   %                 =                    �    �   %                 =                    �    �   %                 =                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�{     �   �   �   �      !                            state�   �   �   �                                  �   �   �   �    5��    �                      G                     �    �                      G                     �    �                     G                    �    �                    c                     �    �                     d                    �    �                     �                     �    �                     �                     �    �                    �                    �    �   '                  �                     �    �   &                  �                     �    �   %                  �                     �    �   $                  �                     �    �   #                  �                     �    �   "                  �                     �    �   !                  �                     �    �                      �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                      �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   �   ,    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    fĶ     �   �   �   �      >                            serial_o <= bit(unsigned(PARITY));5��    �   ,                  j                     5�_�   �   �           �   �   8    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    fĻ     �   �   �   �      A                            serial_o <= bit(to_unsigned(PARITY));5��    �   8                  v                     5�_�   �              �   �   8    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    fĽ     �   �   �   �      D                            serial_o <= bit(to_unsigned(1, PARITY));5��    �   8                  v                     5�_�   �                �   >    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    fĿ     �   �   �   �      A                            serial_o <= bit(to_unsigned(PARITY));5��    �   >                  |                     5�_�                �   +    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    fŵ     �   �   �   �      D                            serial_o <= bit(to_unsigned(PARITY, 1));5��    �   +                  i                     �    �   .                  l                     �    �   -                  k                     �    �   ,                  j                     �    �   +                  i                     �    �   *                  h                     �    �   )                  g                     �    �   (              
   f             
       �    �   (       
          f      
              �    �   (              
   f             
       5�_�    	             ;        ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f�     �   :   <   �    5��    :                      8                     �    :                      8                     �    :                      8                     5�_�    
        	   ;        ����                                                                                                                                                                                                                                                                                                                g   '       z   1       |          V   B    f�     �   ;   G   �          �   <   =   �    �   ;   =   �    5��    ;                      9                     �    ;                      9                     �    ;              
      =              >      5�_�  	            
   =        ����                                                                                                                                                                                                                                                                                                                r   '       =           F                   f�     �   =   G   �   	       if input_int = 0 then           return '0';       elsif input_int = 1 then           return '1';       else   <        -- Handle the case when the input is neither 0 nor 1   7        return '0';  -- or any default value you prefer       end if;   end function int_to_bit;�   <   >   �      begin5��    <                      t                     �    =                      ~                     �    >                      �                     �    ?                      �                     �    @                      �                     �    A                      �                     �    B                      �                     �    C                      ;                     �    D                      w                     �    E                      �                     5�_�  
               C        ����                                                                                                                                                                                                                                                                                                                r   '       =           F                   f�(     �   B   C          @            -- Handle the case when the input is neither 0 nor 15��    B                      �      A               5�_�                 C       ����                                                                                                                                                                                                                                                                                                                q   '       =           E                   f�+     �   B   D   �      ;            return '0';  -- or any default value you prefer5��    B          $                 $               5�_�                 <        ����                                                                                                                                                                                                                                                                                                                q   '       <          <          V       f�K     �   ;   <          :    function int_to_bit(input_int : integer) return bit is   	    begin           if input_int = 0 then               return '0';            elsif input_int = 1 then               return '1';           else               return '0';           end if;       end function int_to_bit;    5��    ;                      9                    5�_�                 J       ����                                                                                                                                                                                                                                                                                                                f   '       <          <          V       f�P     �   J   L   �          �   J   L   �    5��    J                      *                     �    J                     .                     �    J                    A                    �    J                    H                    �    J                      J                     �    J                    I                    �    J   $                  N                     �    J   #                  M                     �    J   "                  L                     �    J   !                  K                     �    J                      J                     �    J                     I                     �    J                 
   H             
       �    J          
          H      
              �    J                 
   H             
       5�_�                 K   (    ����                                                                                                                                                                                                                                                                                                                g   '       <          <          V       f�c     �   J   L   �      (    signal par: bit_vector := bit_vector5��    J   (                  R                     5�_�                 K   )    ����                                                                                                                                                                                                                                                                                                                g   '       <          <          V       f�d     �   J   L   �      *    signal par: bit_vector := bit_vector()5��    J   )                  S                     �    J   )                 S                    �    J   )                 S                    �    J   )                 S                    �    J   )                 S                    5�_�                 K   2    ����                                                                                                                                                                                                                                                                                                                g   '       K   2       K   2       v   2    f�h     �   J   L   �      >    signal par: bit_vector := bit_vector(unsigned(7 downto 0))5��    J   2       
          \      
              �    J   3                  ]                     �    J   2                 \                    �    J   2                 \                    �    J   2              	   \             	       5�_�                 K   )    ����                                                                                                                                                                                                                                                                                                                g   '       K   2       K   2       v   2    f�p     �   J   L   �      =    signal par: bit_vector := bit_vector(unsigned(PARITY, 1))5��    J   )                  S                     5�_�                 K   @    ����                                                                                                                                                                                                                                                                                                                g   '       K   2       K   2       v   2    f�u     �   J   L   �      @    signal par: bit_vector := bit_vector(to_unsigned(PARITY, 1))5��    J   @                  j                     5�_�                 �   (    ����                                                                                                                                                                                                                                                                                                                g   '       K   2       K   2       v   2    fƀ     �   �   �   �      K                            serial_o <= bit_vector(to_unsigned(PARITY, 1));5��    �   (       "          �      "              �    �   *                 �                    5�_�                 �   +    ����                                                                                                                                                                                                                                                                                                                g   '       K   2       K   2       v   2    fƂ     �   �   �   �      ,                            serial_o <= par;5��    �   +                  �                     5�_�                 �   ,    ����                                                                                                                                                                                                                                                                                                                g   '       K   2       K   2       v   2    fƂ     �   �   �   �      .                            serial_o <= par();5��    �   ,                  �                     5�_�                 �   /    ����                                                                                                                                                                                                                                                                                                                g   '       K   2       K   2       v   2    fƞ     �   �   �   �      /                            serial_o <= par(0);5��    �   /                  �                     �    �   3              
   �             
       5�_�                 �   ,    ����                                                                                                                                                                                                                                                                                                                g   '       K   2       K   2       v   2    fƥ    �   �   �   �      ,                            serial_o <= '1';5��    �   ,                                       5�_�                 K       ����                                                                                                                                                                                                                                                                                                                g   '       K   2       K   2       v   2    f�*     �   J   L   �      A    signal par: bit_vector := bit_vector(to_unsigned(PARITY, 1));5��    J                     D                     5�_�                 K       ����                                                                                                                                                                                                                                                                                                                g   '       K   2       K   2       v   2    f�*     �   J   L   �      C    signal par: bit_vector() := bit_vector(to_unsigned(PARITY, 1));5��    J                     E                     5�_�    Z             K       ����                                                                                                                                                                                                                                                                                                                g   '       K   2       K   2       v   2    f�.    �   J   L   �      D    signal par: bit_vector(0) := bit_vector(to_unsigned(PARITY, 1));5��    J                 
   E             
       5�_�    [        Z   �   (    ����                                                                                                                                                                                                                                                                                                                g   '       �   (       �   *       v   *    f�0     �   �   �   �      =                            serial_o <= par(0); -- parity bit�   �   �   �    5��    �   (              "   �             "       5�_�  Z  \          [   K   I    ����                                                                                                                                                                                                                                                                                                                g   '       �   (       �   I       v   *    f�9     �   J   K          M    signal par: bit_vector(0 downto 0) := bit_vector(to_unsigned(PARITY, 1));5��    J                      *      N               5�_�  [  ]          \   ^        ����                                                                                                                                                                                                                                                                                                                f   '       b          h          V       fϏ     �   ^   f   �    �   ^   _   �    5��    ^                      �	              �       5�_�  \  ^          ]   _       ����                                                                                                                                                                                                                                                                                                                m   '       _          e                 fϓ     �   ^   `   �      '                        tx_done <= '1';5��    ^                     �	                     5�_�  ]  _          ^   _       ����                                                                                                                                                                                                                                                                                                                m   '       _          e                 fϕ     �   ^   `   �      #                    tx_done <= '1';5��    ^                     �	                     5�_�  ^  `          _   `       ����                                                                                                                                                                                                                                                                                                                m   '       `          e                 fϛ     �   _   a   �      (                        serial_o <= '1';5��    _                     �	                     5�_�  _  a          `   b       ����                                                                                                                                                                                                                                                                                                                m   '       `          e                 fϝ     �   a   c   �      "                        -- Control5��    a                     �	                     5�_�  `  b          a   c       ����                                                                                                                                                                                                                                                                                                                m   '       `          e                 fϞ     �   b   d   �      ,                        start_signal <= '0';5��    b                    �	                    5�_�  a  c          b   d       ����                                                                                                                                                                                                                                                                                                                m   '       `          e                 fϠ     �   c   e   �      *                        start_stop <= '0';5��    c                     
                     5�_�  b  d          c   d       ����                                                                                                                                                                                                                                                                                                                m   '       `          e                 fϣ     �   c   e   �      +                        Istart_stop <= '0';5��    c          	           
      	               5�_�  c  e          d   e       ����                                                                                                                                                                                                                                                                                                                m   '       `          e                 fϥ   	 �   d   f   �      0                        word <= (others => '0');5��    d                     5
                     5�_�  d  f          e   i        ����                                                                                                                                                                                                                                                                                                                m   '       i          o          V       f��     �   h   i          '                        tx_done <= '1';   (                        serial_o <= '1';       "                        -- Control   ,                        start_signal <= '0';   *                        start_stop <= '0';   0                        word <= (others => '0');5��    h                      �
      �               5�_�  e  g          f   �        ����                                                                                                                                                                                                                                                                                                                    '       i          i          V       f��     �   �   �   �    �   �   �   �    5��    �                      �              �       5�_�  f  h          g   �       ����                                                                                                                                                                                                                                                                                                                    '       �          �                 f��     �   �   �   �      (                        serial_o <= '1';       "                        -- Control   ,                        start_signal <= '0';   *                        start_stop <= '0';   0                        word <= (others => '0');�   �   �   �      '                        tx_done <= '1';5��    �                     �                     �    �                     �                     �    �                     �                     �    �                     #                     �    �                     T                     �    �                     �                     5�_�  g  i          h   i        ����                                                                                                                                                                                                                                                                                                                    '       �          �                 f��     �   h   i           5��    h                      �
                     5�_�  h  j          i   m        ����                                                                                                                                                                                                                                                                                                                    '       m          r          V       f��     �   l   m          '                        tx_done <= '0';   (                        serial_o <= '0';       "                        -- Control   ,                        start_signal <= '1';   %                        word <= data;5��    l                      >      �               5�_�  i  k          j   j        ����                                                                                                                                                                                                                                                                                                                    '       m          m          V       f��     �   j   q   �    �   j   k   �    5��    j                      �
              �       5�_�  j  l          k   k       ����                                                                                                                                                                                                                                                                                                                    '       k          p                 f�      �   k   q   �      (                        serial_o <= '0';       "                        -- Control   ,                        start_signal <= '1';   %                        word <= data;�   j   l   �      '                        tx_done <= '0';5��    j                                          �    k                     =                     �    m                     k                     �    n                     �                     �    o                     �                     5�_�  k  m          l   s        ����                                                                                                                                                                                                                                                                                                                    '       k          p                 f�     �   r   s           5��    r                                           5�_�  l  n          m   u       ����                                                                                                                                                                                                                                                                                                                    '       u          u          V       f�     �   t   u          C                        serial_o <= word(WIDTH-1-signal_bits_sent);5��    t                      h      D               5�_�  m  o          n   s        ����                                                                                                                                                                                                                                                                                                                    '       u          u          V       f�     �   s   u   �    �   s   t   �    5��    s                      D              D       5�_�  n  p          o   x       ����                                                                                                                                                                                                                                                                                                                    '       v          v          V       f�     �   x   z   �    �   x   y   �    5��    x                                    D       5�_�  o  q          p   y       ����                                                                                                                                                                                                                                                                                                                    '       v          v          V       f�)     �   x   z   �      C                        serial_o <= word(WIDTH-1-signal_bits_sent);5��    x                     %                     5�_�  p  s          q           ����                                                                                                                                                                                                                                                                                                                    '                 �          V       f�?     �   ~                                     -- Data   2                        if stop_bits_sent = 0 then   \                            serial_o <= bit_vector(to_unsigned(PARITY, 1))(0); -- parity bit                           else   9                            serial_o <= '1'; -- stop bits                           end if;5��    ~                            '              5�_�  q  t  r      s   |        ����                                                                                                                                                                                                                                                                                                                    '                           V       f�X     �   |   �   �    �   |   }   �    5��    |                      �              '      5�_�  s  u          t   �       ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       f�f     �   �   �   �    �   �   �   �    5��    �                      �              '      5�_�  t  v          u   �       ����                                                                                                                                                                                                                                                                                                                    '       �          �                 f�j     �   �   �   �      2                        if stop_bits_sent = 0 then   \                            serial_o <= bit_vector(to_unsigned(PARITY, 1))(0); -- parity bit                           else   9                            serial_o <= '1'; -- stop bits                           end if;�   �   �   �                              -- Data5��    �                     �                     �    �                     �                     �    �                                          �    �                     p                     �    �                     �                     �    �                     �                     5�_�  u  w          v   }       ����                                                                                                                                                                                                                                                                                                                    '       �          }                 f�o     �   }   �   �      2                        if stop_bits_sent = 0 then   \                            serial_o <= bit_vector(to_unsigned(PARITY, 1))(0); -- parity bit                           else   9                            serial_o <= '1'; -- stop bits                           end if;�   |   ~   �                              -- Data5��    |                     �                     �    }                                          �    ~                     C                     �                         �                     �    �                     �                     �    �                                          5�_�  v  x          w   �        ����                                                                                                                                                                                                                                                                                                                    '       �          }                 f�{     �   �   �           5��    �                      T                     5�_�  w  y          x   v        ����                                                                                                                                                                                                                                                                                                                    '       �          }                 fЁ   
 �   u   v           5��    u                      �                     5�_�  x  z          y   ~        ����                                                                                                                                                                                                                                                                                                                    '       �   ,       �   M       v   M    fШ     �   �   �          `                                serial_o <= bit_vector(to_unsigned(PARITY, 1))(0); -- parity bit�   }      �      `                                serial_o <= bit_vector(to_unsigned(PARITY, 1))(0); -- parity bit5��    }   ,       "          V      "              �    �   ,       "                "              5�_�  y  {          z   K       ����                                                                                                                                                                                                                                                                                                                    '       �   ,       �   M       v   M    fЯ     �   J   L   �          �   J   L   �    5��    J                      *                     �    J                     .                     �    J                     1                     �    J                    0                    �    J                     <                     �    J                     ;                     �    J                 
   :             
       �    J                     C                     �    J                     B                     �    J                     A                     �    J                     @                     �    J                     ?                     �    J                     >                     �    J                     =                     �    J                     <                     �    J                     ;                     �    J                 
   :             
       �    J          
          :      
              �    J                 
   :             
       5�_�  z  |          {   K       ����                                                                                                                                                                                                                                                                                                                    '       �   ,       �   M       v   M    fж     �   J   L   �          signal par: bit_vector5��    J                     D                     5�_�  {  }          |   K       ����                                                                                                                                                                                                                                                                                                                    '       �   ,       �   M       v   M    fж     �   J   L   �          signal par: bit_vector()5��    J                     E                     �    J                    E                    �    J                    G                    �    J                    G                    �    J                    G                    5�_�  |  �          }   K   &    ����                                                                                                                                                                                                                                                                                                                    '       �   ,       �   M       v   M    fк    �   J   L   �      &    signal par: bit_vector(0 downto 0)�   K   L   �    5��    J   &                  P                     �    J   &              '   P             '       5�_�  }  �  ~      �   u   0    ����                                                                                                                                                                                                                                                                                                                    '       u   0       u   )       v   )    f�1     �   t   v   �      C                        serial_o <= word(WIDTH-1-signal_bits_sent);5��    t   0                 �                    5�_�  �  �          �   y   4    ����                                                                                                                                                                                                                                                                                                                    '       u   0       u   )       v   )    f�5    �   x   z   �      G                            serial_o <= word(WIDTH-1-signal_bits_sent);5��    x   4                 �                    5�_�  �  �          �   y   2    ����                                                                                                                                                                                                                                                                                                                    '       u   0       u   )       v   )    f�K     �   x   z   �      G                            serial_o <= word(WIDTH-1+signal_bits_sent);5��    x   2                  �                     5�_�  �  �          �   y   2    ����                                                                                                                                                                                                                                                                                                                    '       u   0       u   )       v   )    f�K     �   x   z   �      F                            serial_o <= word(WIDTH1+signal_bits_sent);5��    x   2                  �                     5�_�  �  �          �   u   .    ����                                                                                                                                                                                                                                                                                                                    '       u   0       u   )       v   )    f�N     �   t   v   �      C                        serial_o <= word(WIDTH-1+signal_bits_sent);5��    t   .                  �                     5�_�  �  �          �   u   .    ����                                                                                                                                                                                                                                                                                                                    '       u   0       u   )       v   )    f�N    �   t   v   �      B                        serial_o <= word(WIDTH1+signal_bits_sent);5��    t   .                  �                     5�_�  �  �          �   u   )    ����                                                                                                                                                                                                                                                                                                                    '       u   0       u   )       v   )    f�[     �   t   v   �      A                        serial_o <= word(WIDTH+signal_bits_sent);5��    t   )                  �                     5�_�  �  �          �   u   :    ����                                                                                                                                                                                                                                                                                                                    '       u   0       u   )       v   )    f�]     �   t   v   �      <                        serial_o <= word(+signal_bits_sent);5��    t   :                  �                     5�_�  �  �          �   u   :    ����                                                                                                                                                                                                                                                                                                                    '       u   0       u   )       v   )    f�^     �   t   v   �      =                        serial_o <= word(+signal_bits_sent-);�   u   v   �    5��    t   ;                  �                     5�_�  �  �          �   u   )    ����                                                                                                                                                                                                                                                                                                                    '       u   0       u   )       v   )    f�a     �   t   v   �      B                        serial_o <= word(+signal_bits_sent-WIDTH);5��    t   )                  �                     5�_�  �  �          �   y   -    ����                                                                                                                                                                                                                                                                                                                    '       y   -       y   B       v   B    f�f    �   x   z   �      E                            serial_o <= word(WIDTH+signal_bits_sent);�   y   z   �    5��    x   -                 �                    5�_�  �  �          �   y   =    ����                                                                                                                                                                                                                                                                                                                    '       y   -       y   B       v   B    fт     �   x   z   �      E                            serial_o <= word(signal_bits_sent-WIDTH);5��    x   =                  �                     5�_�  �  �          �   y   =    ����                                                                                                                                                                                                                                                                                                                    '       y   -       y   B       v   B    fу     �   x   z   �      D                            serial_o <= word(signal_bits_sentWIDTH);5��    x   =                  �                     5�_�  �  �          �   u   9    ����                                                                                                                                                                                                                                                                                                                    '       y   -       y   B       v   B    fх     �   t   v   �      A                        serial_o <= word(signal_bits_sent-WIDTH);5��    t   9                  �                     5�_�  �  �          �   u   9    ����                                                                                                                                                                                                                                                                                                                    '       y   -       y   B       v   B    fц    �   t   v   �      @                        serial_o <= word(signal_bits_sentWIDTH);5��    t   9                  �                     5�_�  �  �          �   i       ����                                                                                                                                                                                                                                                                                                                    '       y   -       y   B       v   B    f��     �   h   j   �    5��    h                      �
                     �    h                      �
                     5�_�  �  �          �   s       ����                                                                                                                                                                                                                                                                                                                    '       z   -       z   B       v   B    f��     �   s   u   �    5��    s                      D                     �    s                      D                     5�_�  �  �          �   w       ����                                                                                                                                                                                                                                                                                                                    '       {   -       {   B       v   B    f��     �   w   y   �    5��    w                      �                     �    w                      �                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   B       v   B    f��    �   �   �   �    5��    �                      P                     �    �                     P                    �    �                      P                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   B       v   B    f��    �         �      B            if (counter > 0) or (start = '1' and counter = 0) then5��                      	   �              	       �       #                  �                     �       "                  �                     �       !                  �                     �                         �                    �                         �                    �                         �                    �       +                  �                     �       *                 �                    �       *                 �                    �       *                 �                    �       4                  �                     �       3                  �                     5�_�  �  �          �      3    ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   B       v   B    f�    �         �      Z            if (counter > 0 and counter < MAX_COUNT) or (start = '1' and counter = 0) then5��       3                  �                     5�_�  �  �          �   �   ,    ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   B       v   B    f��    �   �   �   �      A                                serial_o <= par(0); -- parity bit5��    �   ,                  v                     5�_�  �  �  �      �   q   /    ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   B       v   B    f��     �   p   q          0                            start_signal <= '1';5��    p                      �      1               5�_�  �  �          �   t   #    ����                                                                                                                                                                                                                                                                                                                    '       {   -       {   B       v   B    f��     �   t   v   �    �   t   u   �    5��    t                      S              1       5�_�  �  �          �   u       ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   B       v   B    f��    �   t   v   �      0                            start_signal <= '1';5��    t                     k                     5�_�  �  �  �      �   z       ����                                                                                                                                                                                                                                                                                                                    '       z   +       z          v       f�0     �   y   {   �      1                        if done_signal = '0' then5��    y                    &                    �    y                     )                     �    y                     (                     �    y                     '                     �    y                    &                    �    y   *                  5                     �    y   )                  4                     �    y   (                  3                     �    y   '                  2                     �    y   &                  1                     �    y   %                  0                     �    y   $                  /                     �    y   #                  .                     �    y   "                  -                     �    y   !                  ,                     �    y                      +                     �    y                     *                     �    y                     )                     �    y                     (                     �    y                     '                     �    y                    &                    �    y                    &                    �    y                    &                    5�_�  �  �          �   z   .    ����                                                                                                                                                                                                                                                                                                                    '       z   +       z          v       f�8     �   y   {   �      3                        if signal_bits_sent <  then5��    y   .                  9                     5�_�  �  �          �   z   /    ����                                                                                                                                                                                                                                                                                                                    '       z   +       z          v       f�9     �   y   {   �      5                        if signal_bits_sent < () then5��    y   /                  :                     �    y   /                 :                    �    y   /                 :                    �    y   /                 :                    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f�P     �   �   �   �      /                        if done_stop = '0' then5��    �                    �                    �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �   (                  �                     �    �   '                  �                     �    �   &                  �                     �    �   %                  �                     �    �   $                  �                     �    �   #                  �                     �    �   "                  �                     �    �   !                  �                     �    �                      �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    �    �   /                  �                     �    �   .                  �                     �    �   -                  �                     �    �   ,                 �                    �    �   /                  �                     �    �   .                  �                     �    �   -                  �                     �    �   ,                 �                    �    �   9                  �                     �    �   8                  �                     �    �   7                  �                     �    �   6                  �                     �    �   4                  �                     �    �   3                  �                     �    �   2                  �                     �    �   1                  �                     �    �   0                  �                     �    �   /                  �                     �    �   .                  �                     �    �   -                  �                     �    �   ,                 �                    �    �   ,              	   �             	       �    �   ,       	       	   �      	       	       �    �   ,       	          �      	              �    �   ,              	   �             	       5�_�  �  �          �   z   6    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f�l     �   y   {   �      <                        if signal_bits_sent < (WIDTH-1) then5��    y   6                  A                     5�_�  �  �          �   z   .    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f�n     �   y   {   �      ;                        if signal_bits_sent < (WIDTH-1 then5��    y   .                  9                     5�_�  �  �          �   z   ,    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f�o    �   y   {   �      :                        if signal_bits_sent < WIDTH-1 then5��    y   ,                 7                    5�_�  �  �          �   �   ,    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �   �      A                                serial_o <= par(0); -- parity bit5��    �   ,                  �                     5�_�  �  �          �   �   /    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �          6                            if stop_bits_sent = 0 then5��    �                      S      7               5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �                                       else5��    �                      �      !               5�_�  �  �          �   �   /    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �          =                                serial_o <= '1'; -- stop bits5��    �                      �      >               5�_�  �  �          �   �   "    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �          #                            end if;5��    �                      �      $               5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �   �      E                                serial_o <= not par(0); -- parity bit5��    �                     o                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �          E                                serial_o <= not par(0); -- parity bit5��    �                      �      F               5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �          6                            if stop_bits_sent = 0 then5��    �                      i      7               5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �                                       else5��    �                      i      !               5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �          #                            end if;5��    �                      �      $               5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��    �   �   �   �      =                                serial_o <= '1'; -- stop bits5��    �                     �                     5�_�  �  �          �   z   -    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   y   {   �      :                        if signal_bits_sent = WIDTH-1 then5��    y   ,                 7                    5�_�  �  �          �   z   .    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   y   {   �      :                        if signal_bits_sent < WIDTH-1 then5��    y   .                  9                     5�_�  �  �          �   z   6    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   y   {   �      ;                        if signal_bits_sent < (WIDTH-1 then5��    y   6                  A                     5�_�  �  �  �      �   �   ,    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �   �      :                        if stop_bits_sent = STOP_BITS then5��    �   ,                  	                     5�_�  �  �          �   �   -    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �   �      ;                        if stop_bits_sent = (STOP_BITS then5��    �                     �      <       =       5�_�  �  �          �   �   6    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �   �      <                        if stop_bits_sent = (STOP_BITS) then5��    �   6                                       5�_�  �  �          �   �   6    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �   �      >                        if stop_bits_sent = (STOP_BITS-1) then5��    �   6                                       5�_�  �  �          �   �   6    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �   �      =                        if stop_bits_sent = (STOP_BITS1) then5��    �   6                                       5�_�  �  �          �   �   +    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��    �   �   �   �      <                        if stop_bits_sent = (STOP_BITS) then5��    �   *                                     5�_�  �  �          �   |   $    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f�s     �   |   ~   �    �   |   }   �    5��    |                      �              -       5�_�  �  �          �   }       ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f�t     �   |   ~   �      ,                        start_signal <= '1';5��    |                     �                     5�_�  �  �          �   }   -    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f�w     �   |   ~   �      0                            start_signal <= '1';5��    |   -                 �                    5�_�  �  �          �   �   -    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �   �    �   �   �   �    5��    �                      z              /       5�_�  �  �          �   �   +    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��    �   �   �   �      .                            start_stop <= '1';5��    �   +                 �                    5�_�  �  �          �   w   )    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   v   x   �      ;                        serial_o <= word(signal_bits_sent);5��    v   )                  �                     �    v   *                  �                     �    v   )                 �                    �    v   )                 �                    �    v   )                 �                    5�_�  �  �          �   |   -    ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   <       v   <    f��    �   {   }   �      ?                            serial_o <= word(signal_bits_sent);�   |   }   �    5��    {   -                 �                    5�_�  �  �          �   w   )    ����                                                                                                                                                                                                                                                                                                                    '       w   )       w   0       v   0    f�?     �   v   x   �      C                        serial_o <= word(WIDTH-1-signal_bits_sent);5��    v   )                  �                     5�_�  �  �          �   |   -    ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   4       v   4    f�E     �   {   }   �      G                            serial_o <= word(WIDTH-1-signal_bits_sent);5��    {   -                  �                     5�_�  �  �          �   u   +    ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   4       v   4    f��     �   t   u          ,                        start_signal <= '1';5��    t                      S      -               5�_�  �  �  �      �   p   %    ����                                                                                                                                                                                                                                                                                                                    '       {   -       {   4       v   4    f��     �   p   r   �    �   p   q   �    5��    p                      �              -       5�_�  �  �          �   q       ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   4       v   4    f��     �   p   r   �      ,                        start_signal <= '1';5��    p                     �                     5�_�  �  �          �   }       ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   4       v   4    f��     �   |   }          0                            start_signal <= '0';5��    |                      �      1               5�_�  �  �          �   w       ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   4       v   4    f��     �   w   y   �    �   w   x   �    5��    w                      �              1       5�_�  �  �          �   x       ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f��    �   w   y   �      0                            start_signal <= '0';5��    w                                          5�_�  �  �          �   {   4    ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f�6     �   z   |   �      <                        if signal_bits_sent < (WIDTH-1) then5��    z   4                  p                     5�_�  �  �          �   {   4    ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f�6     �   z   |   �      ;                        if signal_bits_sent < (WIDTH1) then5��    z   4                  p                     5�_�  �  �          �   {   4    ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f�7     �   z   |   �      :                        if signal_bits_sent < (WIDTH) then5��    z   4                  p                     5�_�  �  �          �   {   .    ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f�8    �   z   |   �      9                        if signal_bits_sent < (WIDTH then5��    z   .                  j                     5�_�  �  �          �   T       ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f��    �   S   U   �              generic map(WIDTH)5��    S                     f                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f�=     �   �   �   �                                  �   �   �   �    5��    �                      �                     �    �                     �                     �    �   !                  �                     �    �                      �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�  �  �          �   �   0    ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f�C     �   �   �   �      0                            if stop_bits_sent = 5��    �   0                  �                     5�_�  �  �          �   �   1    ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f�E     �   �   �   �      2                            if stop_bits_sent = ()5��    �   1                  �                     �    �   1              	   �             	       �    �   1       	       	   �      	       	       �    �   1       	          �      	              �    �   1                 �                    5�_�  �  �          �   �   =    ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f�N     �   �   �   �      =                            if stop_bits_sent = (STOP_BITS-1)5��    �   =                  �                     �    �   >                 �                    �    �   >                 �                    �    �   >                 �                    �    �   B                 �                     �    �                  (   �             (       �    �   '                                       �    �   &                                     5�_�  �  �          �   �   "    ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f�X     �   �   �   �      '                                enf if;5��    �   "                                     5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f�X     �   �   �   �      '                                end if;5��    �                                          5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f�[     �   �   �          +                            tx_done <= '1';5��    �                      �      ,               5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f�^     �   �   �   �    �   �   �   �    5��    �                      �              ,       5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                    '       }   -       }   4       v   4    f�`    �   �   �   �      +                            tx_done <= '1';5��    �                                          5�_�  �  �  �      �   �        ����                                                                                                                                                                                                                                                                                                                    '       k          s          V       f@�     �   �   �   �    �   �   �   �    5��    �               	       �              W      5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                    '       �          �                 f@�     �   �   �   �      .                            state <= starting;   +                            tx_done <= '0';   ,                            serial_o <= '0';       &                            -- Control   0                            start_signal <= '1';   )                            word <= data;                           end if;�   �   �   �      +                        if tx_go = '1' then5��    �                     �                     �    �                                          �    �                     4                     �    �                     d                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     $                     5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       f@�     �   �   �          *                            state <= idle;   ,                            serial_o <= '1';       &                            -- Control   0                            start_signal <= '0';   .                            start_stop <= '0';   4                            word <= (others => '0');�   �   �   �      *                            state <= idle;   ,                            serial_o <= '1';       &                            -- Control   0                            start_signal <= '0';   .                            start_stop <= '0';   4                            word <= (others => '0');�   �   �   �    5��   �              �       0                  �    �                                           �    �                      ;                     �    �                      �                     �    �                      �                     �    �                      �                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       f@�     �   �   �   �                                       �   �   �   �    5��    �                                    !       �    �                      ,                     �    �                                           5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       f@�     �   E   H   �          �   E   G   �    5��    E                      �                     �    E                      �                     �    E                     �                     �    F                     �                     �    F                    �                    5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       fA     �   G   P   �          �   H   I   �    �   G   I   �    5��    G                      �                     �    G                    �              �       5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       fA     �   F   G              func5��    F                      �      	               5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       fA     �   F   H   �      6    function natural_to_bit(n : natural) return bit is5��    F                    �                    5�_�  �  �          �   G   *    ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       fA@     �   F   H   �      C    function natural_to_bit(data_to_parity : natural) return bit is5��    F   *                  �                     5�_�  �  �          �   G   ,    ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       fAA     �   F   H   �      B    function natural_to_bit(data_to_parity: natural) return bit is5��    F   ,                 �                    �    F   ,              
   �             
       �    F   ,       
          �      
              �    F   ,              
   �             
       5�_�  �  �          �   G   6    ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       fAC     �   F   H   �      E    function natural_to_bit(data_to_parity: bit_vector) return bit is5��    F   6                  �                     5�_�  �  �          �   G   7    ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       fAE     �   F   H   �      G    function natural_to_bit(data_to_parity: bit_vector()) return bit is5��    F   7                  �                     �    F   8                  �                     �    F   7                 �                    �    F   7                 �                    �    F   7                 �                    �    F   ?                 �                    �    F   ?                 �                    �    F   ?                 �                    5�_�  �  �          �   H       ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       fAu     �   H   J   �    5��    H                      �                     �    H                     �                    5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       fA�     �   H   J   �              5��    H                     �                     �    H                 	   �             	       �    H                    �                    �    H   $                                     �    H   $                                     �    H   $                                     �    H   $                                     �    H   $                                     5�_�  �  �          �   I   2    ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       fB     �   H   J   �      2        variable xor_result: bit := data_to_parity5��    H   2                                       5�_�  �  �          �   I   3    ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       fB     �   H   J   �      4        variable xor_result: bit := data_to_parity()5��    H   3                                       5�_�  �  �          �   I   5    ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       fB     �   H   J   �      5        variable xor_result: bit := data_to_parity(0)5��    H   5                                       5�_�  �  �          �   I   5    ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       fB/     �   H   I          6        variable xor_result: bit := data_to_parity(0);5��    H                      �      7               5�_�  �  �          �   H       ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       fB0     �   G   I   �    �   H   I   �    5��    G                      �              7       5�_�  �  �          �   K        ����                                                                                                                                                                                                                                                                                                                    '       J          N          V       fBN     �   I   K   �          	if n = 0 then�   J   K                  	return '0';   	    	else           	return '1';       	end if;5��    J                      4      A               �    I                     &                     �    I                     !                    5�_�  �  �          �   J       ����                                                                                                                                                                                                                                                                                                                    '       J          K          V       fBk     �   I   K   �              for 1 5��    I                     /                     �    I                    2                    �    I                    2                    �    I                    2                    �    I                    2                    �    I                    2                    �    I                    2                    5�_�  �  �          �   J       ����                                                                                                                                                                                                                                                                                                                    '       J          K          V       fBx     �   J   L   �                  xor_result�   I   L   �              for 1 to WIDTH-15��    I                     9                     �    I                    >              	       �    J                     ?                    �    J                 
   K             
       �    J          
          K      
              �    J                    K                    5�_�  �  �          �   J       ����                                                                                                                                                                                                                                                                                                                    '       J          L          V       fB�     �   I   K   �              for 1 to WIDTH-1 loop5��    I                     -                     5�_�  �  �          �   K       ����                                                                                                                                                                                                                                                                                                                    '       J          L          V       fB�     �   J   L   �                  xor_result <= 5��    J                     ^                     �    J                     `                     �    J                     _                     �    J                 
   ^             
       �    J          
          ^      
              �    J                    ^                    �    J   ,                  p                     �    J   +                  o                     �    J   *                  n                     �    J   )                 m                    �    J   ,                  p                     �    J   +                  o                     �    J   *                  n                     �    J   )                 m                    �    J   6                  z                     �    J   5                  y                     �    J   4                  x                     �    J   3                  w                     �    J   2                  v                     �    J   1                  u                     �    J   0                  t                     �    J   /                  s                     �    J   .                  r                     �    J   -                  q                     �    J   ,                  p                     �    J   +                  o                     �    J   *                  n                     �    J   )                 m                    �    J   )                 m                    �    J   )                 m                    5�_�  �  �          �   K   7    ����                                                                                                                                                                                                                                                                                                                    '       J          L          V       fB�     �   J   L   �      7            xor_result <= xor_result xor data_to_parity5��    J   7                  {                     5�_�  �  �          �   K   8    ����                                                                                                                                                                                                                                                                                                                    '       J          L          V       fB�     �   J   L   �      9            xor_result <= xor_result xor data_to_parity()5��    J   8                  |                     5�_�  �  �          �   K   :    ����                                                                                                                                                                                                                                                                                                                    '       J          L          V       fB�     �   J   L   �      :            xor_result <= xor_result xor data_to_parity(i)5��    J   :                  ~                     5�_�  �  �          �   K   :    ����                                                                                                                                                                                                                                                                                                                    '       J          L          V       fB�     �   K   M   �                  �   K   M   �    5��    K                      �                     �    K                     �                     �    K                     �                    �    K                     �                     5�_�  �  �          �   L       ����                                                                                                                                                                                                                                                                                                                    '       J          M          V       fB�     �   L   N   �              �   L   N   �    5��    L                      �              	       �    L                     �                     �    L   
                  �                     �    L   	                  �                     �    L                    �                    �    L                    �                    �    L                 
   �             
       �    L                     �                     �    L                     �                     �    L                    �                    �    L                    �                    �    L                    �                    �    L                     �                     �    L                     �                     �    L                     �                     �    L                 
   �             
       �    L          
          �      
              �    L                 
   �             
       5�_�  �  �          �   M       ����                                                                                                                                                                                                                                                                                                                    '       J          N          V       fB�     �   L   N   �              return xor_result5��    L                     �                     5�_�  �  �          �   K       ����                                                                                                                                                                                                                                                                                                                    '       J          N          V       fC�     �   J   L   �      ;            xor_result <= xor_result xor data_to_parity(i);5��    J                     \                     �    J                    [                    5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                    '       J          N          V       fD     �   F   H   �      W    function natural_to_bit(data_to_parity: bit_vector(WIDTH-1 downto 0)) return bit is5��    F                    �                    �    F                     �                     �    F                     �                     �    F                     �                     �    F                    �                    �    F                     �                     �    F                     �                     �    F                     �                     �    F                    �                    �    F                     �                     �    F                     �                     �    F                     �                     �    F                     �                     �    F                     �                     �    F                     �                     �    F                     �                     �    F                     �                     �    F                     �                     �    F                     �                     �    F                     �                     �    F                     �                     �    F                     �                     �    F                    �                    �    F                    �                    �    F                    �                    5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                    '       J          N          V       fD     �   F   H   �      W    function data_to_parity(data_to_parity: bit_vector(WIDTH-1 downto 0)) return bit is5��    F                    �                    5�_�  �  �          �   H   $    ����                                                                                                                                                                                                                                                                                                                    '       J          N          V       fD     �   G   I   �      6        variable xor_result: bit := data_to_parity(0);5��    G   $                 �                    5�_�  �  �          �   K   )    ����                                                                                                                                                                                                                                                                                                                    '       J          N          V       fD     �   J   L   �      ;            xor_result := xor_result xor data_to_parity(i);5��    J   )                 Y                    5�_�  �  �          �   N       ����                                                                                                                                                                                                                                                                                                                    '       J          N          V       fD      �   M   O   �      	end function natural_to_bit;5��    M                     �                     5�_�  �  �          �   N       ����                                                                                                                                                                                                                                                                                                                    '       J          N          V       fD!     �   M   O   �      	end function ;5��    M                     �                     5�_�  �             �   T       ����                                                                                                                                                                                                                                                                                                                    '       J          N          V       fD'     �   S   T          M    signal par: bit_vector(0 downto 0) := bit_vector(to_unsigned(PARITY, 1));5��    S                      X      N               5�_�  �                �   ,    ����                                                                                                                                                                                                                                                                                                                    '       �   ,       �   1       v   1    fD0     �   �   �   �      A                            serial_o <= not par(0); -- parity bit5��    �   ,                 v                    �    �   /                  y                     �    �   .                  x                     �    �   -                  w                     �    �   ,                 v                    �    �   /                  y                     �    �   .                  x                     �    �   -                  w                     �    �   ,                 v                    �    �   9                  �                     �    �   8                  �                     �    �   7                  �                     �    �   6                  �                     �    �   5                                       �    �   4                  ~                     �    �   3                  }                     �    �   2                  |                     �    �   1                  {                     �    �   0                  z                     �    �   /                  y                     �    �   .                  x                     �    �   -                  w                     �    �   ,                 v                    �    �   ,                 v                    �    �   ,                 v                    5�_�                  �   :    ����                                                                                                                                                                                                                                                                                                                    '       �   ,       �   1       v   1    fD5     �   �   �   �      I                            serial_o <= not data_to_parity; -- parity bit5��    �   :                  �                     5�_�                   �   ;    ����                                                                                                                                                                                                                                                                                                                    '       �   ,       �   1       v   1    fD6   ! �   �   �   �      K                            serial_o <= not data_to_parity(); -- parity bit5��    �   ;                  �                     �    �   ;                 �                    �    �   ;                 �                    �    �   ;                 �                    5�_�  �      �  �  �   �        ����                                                                                                                                                                                                                                                                                                                    '       k          s          V       f@�     �   �   �   �    �   �   �   �   	   +                        if tx_go = '1' then   .                            state <= starting;   +                            tx_done <= '0';   ,                            serial_o <= '0';       &                            -- Control   0                            start_signal <= '1';   )                            word <= data;                           end if;5��    �               	       �              W      5�_�  �      �  �  �   �        ����                                                                                                                                                                                                                                                                                                                    '       k          s          V       f@�     �   �   �   �                                  �   �   �   �                                  if 5��    �                      �                     �    �                     �                     5�_�  �          �  �   s       ����                                                                                                                                                                                                                                                                                                                    '       �          �          V       f�-     �   r   s   �                                  �   r   t   �                              else    5��    r                      @                     �    r                      @                     �    r                     @                    �    r                     \                     �    r                     \                     �    r                    \                     �    s                     ]                    �    s                      ]                     5�_�  �          �  �   n   (    ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   4       v   4    f��     �   n   o   �    �   n   o   �      ,                        start_signal <= '1';5��    n                      �              -       5�_�  �          �  �   �   ,    ����                                                                                                                                                                                                                                                                                                                    '       �   )       �          v       f��     �   �   �   �      C                        if stop_bits_sent = (((((((((STOP_BITS then5��    �   ,               	   	              	       5�_�  �  �      �  �   x        ����                                                                                                                                                                                                                                                                                                                    '       {   -       {   B       v   B    f��     �   w   y        5��    w                      �                     5�_�  �              �   u       ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   B       v   B    f��     �   t   u   �       5��    t                      S                     �    t                      S                     5�_�  �  �      �  �      5    ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   B       v   B    f�7     �         �      Z            if (counter > 0 and counter < MAX_COUNT) or (start = '1' and counter = 0) then5��       4                  �                     �       3                  �                     5�_�  �              �      $    ����                                                                                                                                                                                                                                                                                                                    '       |   -       |   B       v   B    f�?    �         �      '            if counter = MAX_COUNT then5��       !                 ^                    5�_�  }        �  ~   u   )    ����                                                                                                                                                                                                                                                                                                                    '       y   -       y   4       v   4    f�     �   t   v   �      ;                        serial_o <= word(signal_bits_sent);5��    t   )                  �                     5�_�  ~                 y   -    ����                                                                                                                                                                                                                                                                                                                    '       y   -       y   4       v   4    f�    �   x   z   �      ?                            serial_o <= word(signal_bits_sent);5��    x   -                                       5�_�  q          s  r   �        ����                                                                                                                                                                                                                                                                                                                    '                           V       f�A     �   �   �   �    �   �   �   �                              -- Data   2                        if stop_bits_sent = 0 then   \                            serial_o <= bit_vector(to_unsigned(PARITY, 1))(0); -- parity bit                           else   9                            serial_o <= '1'; -- stop bits                           end if;5��    �                      u              '      5�_�          Z     ^        ����                                                                                                                                                                                                                                                                                                                e   '       ^           ^           V        fʚ     �   ]   `        5��    ]                      �	      J               5�_�                 ]        ����                                                                                                                                                                                                                                                                                                                g   '       ]          ^                 fʛ     �   ]   ^   �    �   \   ]   �                  if reset = '1' then   )                state <= idle; -- repouso5��    \                      a	              J       5�_�                 ]       ����                                                                                                                                                                                                                                                                                                                g   '       ]          ^                 fʣ     �   \   ^   �              if reset = '1' then5��    \                     i	                     5�_�                  ^       ����                                                                                                                                                                                                                                                                                                                g   '       ]          ^                 fʤ     �   ]   _   �      %            state <= idle; -- repouso5��    ]                     �	                     5�_�    !              _       ����                                                                                                                                                                                                                                                                                                                g   '       ]          ^                 fʨ     �   ^   `   �      %        elsif rising_edge(clock) then5��    ^                     �	                     5�_�     "          !   `   
    ����                                                                                                                                                                                                                                                                                                                f   '       ]          ^                 fʪ     �   _   a        5��    _                      �	                     5�_�  !  #          "   _       ����                                                                                                                                                                                                                                                                                                                f   '       ]          ^                 fʫ     �   ^   `   �      )            elsif rising_edge(clock) then5��    ^                     �	                     5�_�  "  $          #   �       ����                                                                                                                                                                                                                                                                                                                f   '       ]          ^                 fʸ     �   �   �   �              end process;5��    �                    1                    �    �                     3                     �    �                     2                     �    �                    1                    �    �                    1                    �    �                    1                    5�_�  #  &          $   �       ����                                                                                                                                                                                                                                                                                                                f   '       ]          �                 fʻ     �   �   �   �          end if;5��    �                    B                    5�_�  $  '  %      &   �       ����                                                                                                                                                                                                                                                                                                                f   '       ]          �                 f��     �   �   �        5��    �                      %                     5�_�  &  (          '   �       ����                                                                                                                                                                                                                                                                                                                f   '       ]          �                 f��     �   �   �   �    �   �   �   �              end process;5��    �                      1                     5�_�  '  )          (   �       ����                                                                                                                                                                                                                                                                                                                f   '       ]          �                 f��     �   �   �   �          end process;5��    �                     5                     5�_�  (  *          )   �       ����                                                                                                                                                                                                                                                                                                                f   '       �          _                 f��     �   �   �   �              end if;5��    �                     )                     5�_�  )  +          *   _       ����                                                                                                                                                                                                                                                                                                                f   '       `          �                 f��     �   ^   `   �      %        elsif rising_edge(clock) then5��    ^                     �	                     5�_�  *  ,          +   `       ����                                                                                                                                                                                                                                                                                                                f   '       `          �                 f�     �   _   a   �                  case state is5��    _                     �	                     5�_�  +  -          ,   a       ����                                                                                                                                                                                                                                                                                                                f   '       `          �                 f�     �   `   b   �                      when idle =>5��    `                     �	                     5�_�  ,  .          -   b       ����                                                                                                                                                                                                                                                                                                                f   '       `          �                 f�     �   a   c   �      #                    tx_done <= '1';5��    a                     
                     5�_�  -  0          .   c       ����                                                                                                                                                                                                                                                                                                                f   '       `          �                 f�     �   b   d   �      $                    serial_o <= '1';5��    b                     8
                     5�_�  .  1  /      0   e       ����                                                                                                                                                                                                                                                                                                                f   '       `          �                 f�
     �   d   f   �                          -- Control5��    d                     ^
                     5�_�  0  2          1   f       ����                                                                                                                                                                                                                                                                                                                f   '       g          h                 f�     �   e   g   �      (                    start_signal <= '0';5��    e                     }
                     5�_�  1  3          2   g       ����                                                                                                                                                                                                                                                                                                                f   '       g          h                 f�     �   f   h   �      &                    start_stop <= '0';5��    f                     �
                     5�_�  2  4          3   h       ����                                                                                                                                                                                                                                                                                                                f   '       g          h                 f�     �   g   i   �      ,                    word <= (others => '0');5��    g                     �
                     5�_�  3  5          4   j       ����                                                                                                                                                                                                                                                                                                                f   '       g          h                 f�     �   i   k   �      '                    if tx_go = '1' then5��    i                     �
                     5�_�  4  6          5   k       ����                                                                                                                                                                                                                                                                                                                f   '       g          h                 f�     �   j   l   �      *                        state <= starting;5��    j                     '                     5�_�  5  7          6   l       ����                                                                                                                                                                                                                                                                                                                f   '       g          h                 f�     �   k   m   �                          end if;5��    k                     N                     5�_�  6  8          7   m   $    ����                                                                                                                                                                                                                                                                                                                f   '       g          h                 f�     �   l   n   �      /                    when starting =>-----------5��    l   $                  z                     5�_�  7  9          8   m   $    ����                                                                                                                                                                                                                                                                                                                f   '       g          h                 f�     �   l   n   �      0                    when starting => -----------5��    l   $                  z                     5�_�  8  :          9   �       ����                                                                                                                                                                                                                                                                                                                f   '       g          h                 f�     �   �   �        5��    �                                           5�_�  9  ;          :   m   $    ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�#     �   l   n   �      $                    when starting =>5��    l   $                  z                     5�_�  :  <          ;   m       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�)     �   l   n   �                       when starting =>5��    l                     f                     5�_�  ;  =          <   n       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�+     �   m   o   �      #                    tx_done <= '0';5��    m                     �                     5�_�  <  >          =   o       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�,     �   n   p   �      $                    serial_o <= '0';5��    n                     �                     5�_�  =  ?          >   q       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�<     �   p   r   �                          -- Control5��    p                     �                     5�_�  >  @          ?   r       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�=     �   q   s   �      (                    start_signal <= '1';5��    q                     �                     5�_�  ?  A          @   s       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�>     �   r   t   �      !                    word <= data;5��    r                                          5�_�  @  B          A   u       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�?     �   t   v   �      %                    state <= sending;5��    t                     @                     5�_�  A  C          B   v       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�@     �   u   w   �                      when sending =>5��    u                     b                     5�_�  B  D          C   w       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�A     �   v   x   �      ?                    serial_o <= word(WIDTH-1-signal_bits_sent);5��    v                     �                     5�_�  C  E          D   y       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�B     �   x   z   �      -                    if done_signal = '0' then5��    x                     �                     5�_�  D  F          E   {       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�C     �   z   |   �                          else5��    z                     #                     5�_�  E  G          F   z       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�D     �   y   {   �      )                        state <= sending;5��    y                     �                     5�_�  F  H          G   |       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�G     �   {   }   �      *                        state <= stopping;5��    {                     <                     5�_�  G  I          H   }       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�H     �   |   ~   �      *                        start_stop <= '1';5��    |                     g                     5�_�  H  J          I   ~       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�I     �   }      �                          end if;5��    }                     �                     5�_�  I  K          J          ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�J     �   ~   �   �                       when stopping =>5��    ~                     �                     5�_�  J  L          K   �       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�K     �      �   �                          -- Data5��                         �                     5�_�  K  M          L   �       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�L     �   �   �   �      .                    if stop_bits_sent = 0 then5��    �                     �                     5�_�  L  N          M   �       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�M     �   �   �   �      9                        serial_o <= par(0); -- parity bit5��    �                                          5�_�  M  O          N   �       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�O     �   �   �   �                          else5��    �                     P                     5�_�  N  P          O   �       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�P     �   �   �   �      5                        serial_o <= '1'; -- stop bits5��    �                     m                     5�_�  O  R          P   �       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�Q     �   �   �   �                          end if;5��    �                     �                     5�_�  P  S  Q      R   �       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�T     �   �   �   �      +                    if done_stop = '0' then5��    �                     �                     5�_�  R  T          S   �       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�U     �   �   �   �      *                        state <= stopping;5��    �                     �                     5�_�  S  U          T   �       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�V     �   �   �   �                          else5��    �                                          5�_�  T  V          U   �       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�W     �   �   �   �      &                        state <= idle;5��    �                     0                     5�_�  U  W          V   �       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�X     �   �   �   �                          end if;5��    �                     S                     5�_�  V  X          W   �       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�Y     �   �   �   �                  end case;5��    �                     g                     5�_�  W  Y          X   �       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�Z    �   �   �   �              end if;5��    �                     y                     5�_�  X              Y   [       ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 fͺ    �   Z   \   �      #    process(clock, reset, tx_go) is5��    Z                     R	                     �    Z                     \	                     �    Z                    [	                    �    Z                    [	                    �    Z                    [	                    �    Z                    [	                    �    Z                    [	                    5�_�  P          R  Q   �        ����                                                                                                                                                                                                                                                                                                                f   '       m          �                 f�R     �   �   �   �       �   �   �   �                          end if;5��    �                     �                     5�_�  .          0  /   d        ����                                                                                                                                                                                                                                                                                                                e   '       `          �                 f�     �   c   e   �       �   b   e   �      $                    serial_o <= '1';5��    b   $                  H
                     5�_�  $          &  %   �       ����                                                                                                                                                                                                                                                                                                                f   '       ]          ^                 f��     �   �   �   �              end process5��    �                     8                     5�_�            	     ;        ����                                                                                                                                                                                                                                                                                                                g   '       z   1       |          V   B    f�     �   ;   <   �    �   :   <   �      15��    :                      8                     5�_�                �   ,    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f��     �   �   �   �      9                            serial_o <= bit((PARITY, 1));5��    �   ,                  j                     5�_�                 �   ,    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f��     �   �   �   �      8                            serial_o <= bit(PARITY, 1));5��    �   ,                  j                     5�_�                 �   6    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f��     �   �   �   �      7                            serial_o <= bit(PARITY, 1);5��    �   6                  t                     5�_�                 �   2    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f��     �   �   �   �      5                            serial_o <= bit(PARITY1);5��    �   2                  p                     5�_�                   �   2    ����                                                                                                                                                                                                                                                                                                                f   '       y   1       {          V   B    f��     �   �   �   �      4                            serial_o <= bit(PARITY);5��    �   2                  p                     5�_�   �           �   �   �       ����                                                                                                                                                                                                                                                                                                                f   '       z   1       |          V   B    f��     �   �   �   �                              5��    �          !                 !               5�_�   �           �   �   g   '    ����                                                                                                                                                                                                                                                                                                                f   '       g   '       e   "       V   '    f��     �   g   h   �       5��    g                      �
                     �    g                      �
                     5�_�   �           �   �   f   '    ����                                                                                                                                                                                                                                                                                                                f   '                                        f�\     �   e   h         ?                        start_signal <= '0'; start_stop <= '0';5��    e   ,                W
                    5�_�   �           �   �   N        ����                                                                                                                                                                                                                                                                                                                            \          M          V       f�B     �   M   O   �      %    signal signal_bits_done: natural;�   Q   S          #    signal stop_bits_done: natural;�   W   Y          P        port map(clock, reset, start_signal, finished_signal, signal_bits_done);�   [   ]          J        port map(clock, reset, start_stop, finished_stop, stop_bits_done);5��    M                    }                    �    Q                    �                    �    W   J                                     �    [   D                 
	                    5�_�   �   �       �   �   C       ����                                                                                                                                                                                                                                                                                                                            =          C                 f��     �   B   D        5��    B                            G               5�_�   �   �           �   #        ����                                                                                                                                                                                                                                                                                                                            ;          A                 f��     �   "   %        5��    "                      _                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            :          @                 f��     �   
           5��    
                      �       C               5�_�   �               �   
       ����                                                                                                                                                                                                                                                                                                                            :          @                 f��     �   	      r              done: out bit5��    	                     �                      5�_�   3           5   4   "       ����                                                                                                                                                                                                                                                                                                                            "   &       "   &       v   &    f�O     �   !   #   .      4                case std_logic_vector(7 downto 0) is5��    !                                        �    !                                        �    !                                        �    !                                        �    !                                        5�_�   $           &   %          ����                                                                                                                                                                                                                                                                                                                                                          f�     �               )    type transmiter is (, sending, idle);5��              	           �      	               5�_�                            ����                                                                                                                                                                                                                                                                                                                                                v       f?r     �               �    signal PALAVRA_TRANSMITIR: std_logic_vector (9 downto 0) := "1111111111"; -- Vetor que guardará a palavra a ser enviada via serial     5��                          �                     5��