Vim�UnDo� �(���$N�Rd�%�jT!#�@��C���   P   H        assert count = "000001" report "Did not proceed" severity error;   J        .      .  .  .    f�o     _�                             ����                                                                                                                                                                                                                                                                                                                                                             f ǌ     �                   �               5��                    =                      m      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f ǟ     �         >      end Temporized_Testbench;5��                         i                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f Ǡ     �         >      end ;5��                         h                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f ǡ     �         >      entity Temporized_Testbench is   end;�         >      end;5��                         d                      �                         d                      5�_�      	                    ����                                                                                                                                                                                                                                                                                                                                                V       f ǰ     �         =      #entity Temporized_Testbench is end;5��                        M                     5�_�      
          	          ����                                                                                                                                                                                                                                                                                                                                                V       f Ǹ     �         =      entity count is end;5��                         R                      5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                         .       v   .    f ��     �         =      2architecture Behavioral of Temporized_Testbench is�         =    5��                     
   |              
       5�_�   
                    $    ����                                                                                                                                                                                                                                                                                                                                         $       v   .    f ��     �      	   =      K    constant CLOCK_PERIOD : time := 10 ns;  -- Clock period (e.g., 100 MHz)5��       $                 �                     5�_�                       C    ����                                                                                                                                                                                                                                                                                                                               C          D       v   D    f ��     �      	   =      K    constant CLOCK_PERIOD : time := 20 ns;  -- Clock period (e.g., 100 MHz)5��       C                 �                     5�_�                    
       ����                                                                                                                                                                                                                                                                                                                               C          D       v   D    f ��     �   	      =      3    signal clk : std_logic := '0';  -- Clock signal5��    	          	          �       	              �    	                     �                      �    	                    �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                               C          D       v   D    f ��     �   
      =      5    signal reset : std_logic := '0';  -- Reset signal5��    
          	                	              5�_�                           ����                                                                                                                                                                                                                                                                                                                               C          D       v   D    f ��     �         =      P    signal stimulus : std_logic_vector(3 downto 0) := "0000";  -- Input stimulus5��                     
   J             
       5�_�                       !    ����                                                                                                                                                                                                                                                                                                                               C          D       v   D    f ��     �         =      J    signal stimulus : bit_vector(3 downto 0) := "0000";  -- Input stimulus5��       !                 U                    5�_�                       1    ����                                                                                                                                                                                                                                                                                                                               C          D       v   D    f ��     �         =      J    signal stimulus : bit_vector(5 downto 0) := "0000";  -- Input stimulus5��       1                  e                     5�_�                       1    ����                                                                                                                                                                                                                                                                                                                               C          D       v   D    f ��     �         =      K    signal stimulus : bit_vector(5 downto 0) := "00000";  -- Input stimulus5��       1                  e                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                         (       v   (    f �    �         =      )    DUT_Instance : entity work.DUT_Entity�         =    5��              
          0      
              5�_�                           ����                                                                                                                                                                                                                                                                                                                                         +       v   (    f�     �         =      ,    DUT_Instance : entity work.counter_6bit 5��                                            5�_�                           ����                                                                                                                                                                                                                                                                                                                                         +       v   (    f�     �         =      #    dut : entity work.counter_6bit 5��                                              5�_�                          ����                                                                                                                                                                                                                                                                                                                                         +       v   (    f�     �      	   =    5��                          �                      �                          �                      �                          �                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                         +       v   (    f�     �      
   ?          �      	   >    5��                          �                      �                          �                      �                          �                      �                         �                      �                      	   �               	       5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                         +       v   (    f�     �   	      @    �   	   
   @    5��    	                      �                     5�_�                    	       ����                                                                                                                                                                                                                                                                                                                            &          &   +       v   (    f�     �      	              component5��                          �                      5�_�                    	       ����                                                                                                                                                                                                                                                                                                                            %          %   +       v   (    f��     �      	          <    -- Component declaration for the DUT (Design Under Test)5��                          �       =               5�_�                            ����                                                                                                                                                                                                                                                                                                                            $          $   +       v   (    f��     �                 5��                          �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f��     �      	   E          component somador�      	   E    5��                        �                     5�_�                    
        ����                                                                                                                                                                                                                                                                                                                            
                    V       f��     �   	      B    �   
      B    �   	   
          +            A : in bit_vector(31 downto 0);   +            B : in bit_vector(31 downto 0);   +            S : out bit_vector(31 downto 0)5��    	                      �       �               �    	                      �               �       5�_�                     
       ����                                                                                                                                                                                                                                                                                                                            
                           f��     �   
      E      =        rst : in bit;                          -- Reset input   Q        count : out bit_vector(5 downto 0)       -- 6-bit count output (64 steps)�   	      E      ?        clk : in bit;                            -- Clock input5��    	                     �                      �    
                                           �                         B                     5�_�      !               "       ����                                                                                                                                                                                                                                                                                                                            
                           f��     �   !   "          :    -- Replace DUT_Entity with the name of your DUT entity5��    !                      �      ;               5�_�       "           !   "   	    ����                                                                                                                                                                                                                                                                                                                            
                           f�      �   !   #   D      "    dut: entity work.counter_6bit 5��    !   	                                     �    !                                          �    !                                          �    !   
                                       �    !   	                                     �    !   	                                     �    !   	                                     5�_�   !   #           "   %       ����                                                                                                                                                                                                                                                                                                                            
                           f�     �   $   &   D                  reset => reset,5��    $                    H                    �    $                     I                     �    $                    H                    �    $                    H                    �    $                    H                    5�_�   "   $           #   &       ����                                                                                                                                                                                                                                                                                                                            
                           f�     �   %   '   D                   stimulus => stimulus5��    %                    b                    �    %                     c                     �    %                    b                    �    %                    b                    �    %                    b                    5�_�   #   %           $   '       ����                                                                                                                                                                                                                                                                                                                            
                           f�     �   &   '          (            -- Add other ports as needed5��    &                      t      )               5�_�   $   &           %   *       ����                                                                                                                                                                                                                                                                                                                            
                           f�     �   )   +   C          stimulus_process: process5��    )                     �                     5�_�   %   (           &   8       ����                                                                                                                                                                                                                                                                                                                            
                           f�$     �   7   9   C      !    end process stimulus_process;5��    7                    �                    5�_�   &   )   '       (   0       ����                                                                                                                                                                                                                                                                                                                            
                           f�G     �   0   2   C    5��    0                      �              	       �    0                      �                     5�_�   (   *           )   0       ����                                                                                                                                                                                                                                                                                                                            
                           f�J     �   /   1   D      0        stimulus <= "0001";  -- Example stimulus5��    /                    �                    5�_�   )   +           *   1        ����                                                                                                                                                                                                                                                                                                                            3          2          V       f�P     �   1   4   D    �   1   2   D    5��    1                      �              P       5�_�   *   ,           +   3       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�T     �   2   4   F      0        stimulus <= "0010";  -- Example stimulus5��    2                    �                    5�_�   +   -           ,   3       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�U     �   2   4   F      0        stimulus <= "0000";  -- Example stimulus5��    2                    �                    5�_�   ,   .           -   7       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�Z     �   6   8   F      0        stimulus <= "0100";  -- Example stimulus5��    6                    �                    5�_�   -   /           .   7       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�[     �   6   8   F      0        stimulus <= "0101";  -- Example stimulus5��    6                    �                    5�_�   .   0           /   7       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�\     �   6   8   F      0        stimulus <= "0111";  -- Example stimulus5��    6                    �                    5�_�   /   1           0   9       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�]     �   8   :   F      0        stimulus <= "1000";  -- Example stimulus5��    8                    �                    5�_�   0   2           1   9       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�^     �   8   :   F      0        stimulus <= "1100";  -- Example stimulus5��    8                    �                    5�_�   1   3           2   9       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�_     �   8   :   F      0        stimulus <= "1100";  -- Example stimulus5��    8                    �                    5�_�   2   4           3   0       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�o     �   /   1   F      0        stimulus <= "0000";  -- Example stimulus5��    /                     �                     5�_�   3   5           4   0       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�p     �   /   1   F              stimulus <= "0000";  5��    /                     �                     5�_�   4   6           5   0       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�p     �   /   1   F              stimulus <= "0000"; 5��    /                     �                     5�_�   5   7           6   3       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�{     �   2   4   F      0        stimulus <= "0001";  -- Example stimulus5��    2                     �                     5�_�   6   8           7   5       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�}     �   4   6   F      0        stimulus <= "0010";  -- Example stimulus5��    4                                          5�_�   7   9           8   7       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�     �   6   8   F      0        stimulus <= "0011";  -- Example stimulus5��    6                     G                     5�_�   8   :           9   9       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�     �   8   :   F      0        stimulus <= "0100";  -- Example stimulus5��    8                     �                     5�_�   9   ;           :   A       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�     �   @   B   F      0        wait for 20 ns;  -- Hold reset for 20 ns5��    @                    %                    �    @                     '                     �    @                     &                     �    @                    %                    �    @                     )                     �    @                     (                     �    @                     '                     �    @                     &                     �    @                    %                    �    @                     )                     �    @                     (                     �    @                     '                     �    @                     &                     �    @                    %                    �    @                    %                    �    @                    %                    �    @                    %                    5�_�   :   <           ;   @       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�     �   ?   A   G              �   ?   A   F    5��    ?                      �              	       �    ?                     �                     �    ?                     �                     �    ?   
                  �                     �    ?   	                  �                     �    ?                    �                    �    ?                     �                     �    ?   
                  �                     �    ?   	                  �                     �    ?                    �                    �    ?                     �                     �    ?                     �                     �    ?                     �                     �    ?                     �                     �    ?                     �                     �    ?   
                  �                     �    ?   	                  �                     �    ?                    �                    �    ?                    �                    �    ?                    �                    5�_�   ;   =           <   @       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�     �   ?   A   G              stimulus <= 5��    ?                                          5�_�   <   ?           =   @       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�     �   ?   A   G              stimulus <= ""5��    ?                                          5�_�   =   @   >       ?   C       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�     �   B   D   H              �   B   D   G    5��    B                      g              	       �    B                     o                     �    B                    o                    �    B                    o                    �    B                    o                    �    B                 2   o             2       5�_�   ?   A           @   C       ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�     �   B   D   H      :        assert neg_condition report message severity note;5��    B                    v                    �    B                     w                     �    B                    v                    5�_�   @   B           A   C       ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�     �   B   D   H      5        assert count =  report message severity note;5��    B                     ~                     5�_�   A   C           B   C       ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�     �   B   D   H      7        assert count = "" report message severity note;5��    B                                          5�_�   B   D           C   0       ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�$     �   /   1   H              stimulus <= "0000";5��    /                     �                     5�_�   C   E           D   3       ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�'     �   2   4   H              stimulus <= "0001";5��    2                     �                     5�_�   D   F           E   5       ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�*     �   4   6   H              stimulus <= "0010";5��    4                     
                     5�_�   E   G           F   7       ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�,     �   6   8   H              stimulus <= "0011";5��    6                     G                     5�_�   F   H           G   9       ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�/     �   8   :   H              stimulus <= "0100";5��    8                     �                     5�_�   G   I           H   @       ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�2     �   ?   A   H              stimulus <= "1011"5��    ?                                          5�_�   H   J           I   @       ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�7     �   ?   A   H              stimulus <= "001011"5��    ?                                          5�_�   I   K           J   C       ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�B     �   B   D   H      =        assert count = "000000" report message severity note;5��    B                    �                    �    B                     �                     �    B                     �                     �    B                     �                     �    B                    �                    �    B                     �                     �    B                     �                     �    B                     �                     �    B                    �                    �    B                     �                     �    B                     �                     �    B                     �                     �    B                     �                     �    B                     �                     �    B                     �                     �    B                     �                     �    B                    �                    �    B                    �                    �    B                    �                    5�_�   J   L           K   C   *    ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�L     �   B   D   H      @        assert stimulus = "000000" report message severity note;5��    B   *                  �                     5�_�   K   M           L   C   *    ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�M     �   B   D   H      9        assert stimulus = "000000" report  severity note;5��    B   *                  �                     5�_�   L   N           M   C   +    ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�Y     �   B   D   H      ;        assert stimulus = "000000" report "" severity note;5��    B   +                  �                     �    B   7                  �                     �    B   6                  �                     �    B   5                  �                     �    B   4                  �                     �    B   3                 �                    �    B   3                 �                    �    B   3                 �                    �    B   C                  �                     �    B   D                  �                     �    B   C                  �                     5�_�   M   O           N   C   C    ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�c     �   B   D   H      H        assert stimulus = "000000" report "Did not reset" severity note;5��    B   C                 �                    �    B   E                 �                    5�_�   N   P           O   D   '    ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�     �   D   F   H    �   D   E   H    5��    D                      �              8       5�_�   O   Q           P   E       ����                                                                                                                                                                                                                                                                                                                            C          C          v       f�     �   E   G   J              �   E   G   I    5��    E                                    	       �    E                     '                     �    E   
                  )                     �    E   	                  (                     �    E                    '                    �    E                    '                    �    E                    '                    �    E                 2   '             2       5�_�   P   R           Q   F       ����                                                                                                                                                                                                                                                                                                                            F          F          v       f�     �   E   G   J      :        assert neg_condition report message severity note;5��    E                    .                    �    E                     0                     �    E                     /                     �    E                    .                    �    E                    .                    �    E                    .                    5�_�   Q   S           R   F       ����                                                                                                                                                                                                                                                                                                                            F          F          v       f�     �   E   G   J      8        assert stimulus =  report message severity note;5��    E                     9                     5�_�   R   T           S   F       ����                                                                                                                                                                                                                                                                                                                            F          F          v       f�     �   E   G   J      :        assert stimulus = "" report message severity note;5��    E                     :                     5�_�   S   U           T   F   *    ����                                                                                                                                                                                                                                                                                                                            F   0       F   *       v   *    f�     �   E   G   J      @        assert stimulus = "000001" report message severity note;5��    E   *                  I                     5�_�   T   V           U   F   *    ����                                                                                                                                                                                                                                                                                                                            F   0       F   *       v   *    f�     �   E   G   J      9        assert stimulus = "000001" report  severity note;5��    E   *                  I                     5�_�   U   W           V   F   +    ����                                                                                                                                                                                                                                                                                                                            F   0       F   *       v   *    f�     �   E   G   J      ;        assert stimulus = "000001" report "" severity note;5��    E   +                  J                     �    E   8                  W                     �    E   7                 V                    �    E   E                  d                     �    E   E                  d                     5�_�   V   X           W   F   E    ����                                                                                                                                                                                                                                                                                                                            F   0       F   *       v   *    f�     �   E   G   J      J        assert stimulus = "000001" report "Did not proceed" severity note;5��    E   E                 d                    5�_�   W   Y           X   3       ����                                                                                                                                                                                                                                                                                                                            F   0       F   *       v   *    f��     �   2   4   J              stimulus <= "000001";5��    2                    �                    �    2   
                  �                     �    2   	                  �                     �    2                    �                    �    2                    �                    �    2                    �                    �    2                 2   �             2       5�_�   X   Z           Y   3       ����                                                                                                                                                                                                                                                                                                                            3          3          v       f��     �   2   4   J      :        assert neg_condition report message severity note;5��    2                    �                    �    2                     �                     �    2                     �                     �    2                    �                    �    2                    �                    �    2                    �                    5�_�   Y   [           Z   3       ����                                                                                                                                                                                                                                                                                                                            3          3          v       f��     �   2   4   J      8        assert stimulus =  report message severity note;5��    2                     �                     5�_�   Z   \           [   3       ����                                                                                                                                                                                                                                                                                                                            3          3          v       f��     �   2   4   J      :        assert stimulus = "" report message severity note;5��    2                     �                     �    2                      �                     �    2                     �                     �    2                     �                     �    2                     �                     �    2                     �                     �    2                    �                    �    2                      �                     �    2                     �                     �    2                     �                     �    2                     �                     �    2                     �                     �    2                    �                    �    2                    �                    �    2                    �                    5�_�   [   ]           \   3   *    ����                                                                                                                                                                                                                                                                                                                            3   0       3   *       v   *    f��     �   2   4   J      @        assert stimulus = "000001" report message severity note;5��    2   *                  �                     5�_�   \   ^           ]   3   *    ����                                                                                                                                                                                                                                                                                                                            3   0       3   *       v   *    f��     �   2   4   J      9        assert stimulus = "000001" report  severity note;5��    2   *                  �                     5�_�   ]   _           ^   3   +    ����                                                                                                                                                                                                                                                                                                                            3   0       3   *       v   *    f��     �   2   4   J      ;        assert stimulus = "000001" report "" severity note;5��    2   +               
   �              
       �    2   4                 �                    �    2   :                  �                     �    2   9                  �                     �    2   8                  �                     �    2   7                 �                    �    2   8                 �                    5�_�   ^   `           _   3   J    ����                                                                                                                                                                                                                                                                                                                            3   0       3   *       v   *    f��     �   2   4   J      O        assert stimulus = "000001" report "Did not proceed to 1" severity note;5��    2   J                                     �    2   K                                     5�_�   _   a           `   4       ����                                                                                                                                                                                                                                                                                                                            3   0       3   *       v   *    f��     �   4   6   J    �   4   5   J    5��    4                      (              Q       5�_�   `   b           a   7       ����                                                                                                                                                                                                                                                                                                                            3   0       3   *       v   *    f��     �   7   9   K    �   7   8   K    5��    7                      �              Q       5�_�   a   c           b   :       ����                                                                                                                                                                                                                                                                                                                            3   0       3   *       v   *    f��     �   :   <   L    �   :   ;   L    5��    :                      D              Q       5�_�   b   d           c   6       ����                                                                                                                                                                                                                                                                                                                            3   0       3   *       v   *    f�     �   5   7   M              stimulus <= "000010";5��    5          	           �      	               5�_�   c   e           d   5       ����                                                                                                                                                                                                                                                                                                                            5          5   "       v   "    f�     �   4   6   M      P        assert stimulus = "000001" report "Did not proceed to 1" severity error;�   5   6   M    5��    4          	       	   B      	       	       5�_�   d   f           e   5   #    ����                                                                                                                                                                                                                                                                                                                            5          5   "       v   "    f�
     �   4   6   M      P        assert stimulus =  "000010"report "Did not proceed to 1" severity error;5��    4   #                  K                     5�_�   e   g           f   5       ����                                                                                                                                                                                                                                                                                                                            5          5   "       v   "    f�     �   4   6   M      Q        assert stimulus =  "000010" report "Did not proceed to 1" severity error;5��    4                     A                     5�_�   f   h           g   5       ����                                                                                                                                                                                                                                                                                                                            5          5   "       v   "    f�     �   4   6   M      O        assert stimulus ="000010" report "Did not proceed to 1" severity error;5��    4                     A                     5�_�   g   i           h   6       ����                                                                                                                                                                                                                                                                                                                            5          5   "       v   "    f�     �   5   6                  stimulus <=;5��    5                      y                     5�_�   h   j           i   8       ����                                                                                                                                                                                                                                                                                                                            5          5   "       v   "    f�     �   7   9   L              stimulus <= "000011";5��    7                     �                     5�_�   i   k           j   7       ����                                                                                                                                                                                                                                                                                                                            7          7           v        f�     �   6   8   L      P        assert stimulus = "000001" report "Did not proceed to 1" severity error;�   7   8   L    5��    6                    �                    5�_�   j   l           k   8       ����                                                                                                                                                                                                                                                                                                                            7          7           v        f�     �   7   8                  stimulus <= "";5��    7                      �                     5�_�   k   m           l   :       ����                                                                                                                                                                                                                                                                                                                            7          7           v        f�&     �   9   ;   K              stimulus <= "000100";5��    9                     n                     5�_�   l   n           m   9       ����                                                                                                                                                                                                                                                                                                                            9          9           v        f�(     �   8   :   K      P        assert stimulus = "000001" report "Did not proceed to 1" severity error;�   9   :   K    5��    8                    #                    5�_�   m   o           n   :       ����                                                                                                                                                                                                                                                                                                                            9          9           v        f�)     �   9   :                  stimulus <= "";5��    9                      Y                     5�_�   n   p           o   5   >    ����                                                                                                                                                                                                                                                                                                                            9          9           v        f�0     �   4   6   J      P        assert stimulus = "000010" report "Did not proceed to 1" severity error;5��    4   >                 f                    5�_�   o   q           p   7   >    ����                                                                                                                                                                                                                                                                                                                            9          9           v        f�1     �   6   8   J      P        assert stimulus = "000011" report "Did not proceed to 1" severity error;5��    6   >                 �                    5�_�   p   v           q   9   >    ����                                                                                                                                                                                                                                                                                                                            9          9           v        f�2    �   8   :   J      P        assert stimulus = "000100" report "Did not proceed to 1" severity error;5��    8   >                 F                    5�_�   q   w   r       v   '   	    ����                                                                                                                                                                                                                                                                                                                            9          9           v        f�p     �   '   *   K              �   '   )   J    5��    '                                    	       �    '                                           �    '                                   	       �    (                     �                     �    (                     �                     �    (                     �                     �    (                    �                    5�_�   v   x           w   )       ����                                                                                                                                                                                                                                                                                                                            ;          ;           v        f��     �   (   )              -- Clock5��    (                      �                     5�_�   w   y           x   )        ����                                                                                                                                                                                                                                                                                                                            :          :           v        f��     �   (   )           5��    (                      �                     5�_�   x   z           y           ����                                                                                                                                                                                                                                                                                                                            9          9           v        f��     �         K          �         J    5��                          �                     �                      
   �              
       �                        �                    �                     
   �             
       �                         �                     �                        �                    �                         �                     �                         �                     �                        �                    �       #                  �                     �       "                  �                     �       !                  �                     �                          �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �                          �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    5�_�   y   {           z      %    ����                                                                                                                                                                                                                                                                                                                            :          :           v        f��     �         K      %    clk <= clk after CLOCK_PERIOD / 25��       %                  �                     5�_�   z   |           {          ����                                                                                                                                                                                                                                                                                                                            :          :           v        f��     �         K      &    clk <= clk after CLOCK_PERIOD / 2)5��                         �                     5�_�   {   }           |      '    ����                                                                                                                                                                                                                                                                                                                            :          :           v        f��     �         K      '    clk <= clk after (CLOCK_PERIOD / 2)5��       '                  �                     5�_�   |   ~           }      '    ����                                                                                                                                                                                                                                                                                                                            :          :           v        f��     �                (    clk <= clk after (CLOCK_PERIOD / 2);5��                          �      )               5�_�   }              ~           ����                                                                                                                                                                                                                                                                                                                            9          9           v        f��     �      !   J    �          J    5��                          �              )       5�_�   ~   �                     ����                                                                                                                                                                                                                                                                                                                                                V       f��    �             	       -- Clock generator process       clk_gen_process: process   	    begin   9        while now < 1000 ns loop  -- Simulate for 1000 ns   ,            clk <= not clk;  -- Toggle clock   E            wait for CLOCK_PERIOD / 2;  -- Wait for half clock period           end loop;           wait;        end process clk_gen_process;5��           	               �      4              5�_�      �           �   1        ����                                                                                                                                                                                                                                                                                                                                      B          V       f��     �   1   3   B    �   1   2   B    5��    1                      N                     5�_�   �   �           �   2       ����                                                                                                                                                                                                                                                                                                                                      C          V       f��     �   2   5   D              �   2   4   C    5��    2                      m              	       �    2                      m                     �    2                     m              	       �    3                     u                     �    3                     t                     �    3                     s                     �    3                     r                     �    3                     q                     �    3                     p                     �    3                     o                     �    3                      n                     5�_�   �   �           �   ;        ����                                                                                                                                                                                                                                                                                                                            ;           A           V        f��     �   :   ;                  stimulus <= "001011";   &        reset <= '1';  -- Assert reset   7        wait for CLOCK_PERIOD;  -- Hold reset for 20 ns   I        assert stimulus = "000000" report "Did not reset" severity error;   (        reset <= '0';  -- Deassert reset   7        wait for CLOCK_PERIOD;  -- Hold reset for 20 ns   K        assert stimulus = "000001" report "Did not proceed" severity error;5��    :                      �      t              5�_�   �   �           �   3        ����                                                                                                                                                                                                                                                                                                                            ;           ;           V        f��     �   3   ;   >    �   3   4   >    5��    3                      n              t      5�_�   �   �           �   ?        ����                                                                                                                                                                                                                                                                                                                            ?          C          V       f��     �   >   ?              -- Reset process (optional)       reset_process: process   	    begin           wait;       end process reset_process;5��    >                            r               5�_�   �   �           �   ?        ����                                                                                                                                                                                                                                                                                                                            ?          ?          V       f��     �   >   ?           5��    >                                           5�_�   �   �           �   >        ����                                                                                                                                                                                                                                                                                                                            ?          ?          V       f��    �   =   >           5��    =                                           5�_�   �   �           �   :        ����                                                                                                                                                                                                                                                                                                                            4           :           V        f��    �   3   ;   >              stimulus <= "001011";   &        reset <= '1';  -- Assert reset   7        wait for CLOCK_PERIOD;  -- Hold reset for 20 ns   I        assert stimulus = "000000" report "Did not reset" severity error;   (        reset <= '0';  -- Deassert reset   7        wait for CLOCK_PERIOD;  -- Hold reset for 20 ns   K        assert stimulus = "000001" report "Did not proceed" severity error;5��    3                     n      t      �      5�_�   �   �           �   (        ����                                                                                                                                                                                                                                                                                                                            4           :           V        f��    �   '   )   >              stimulus <= "000000";5��    '                     o             !       5�_�   �   �           �   +   ?    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f�>     �   *   ,   >      P        assert stimulus = "000001" report "Did not proceed to 1" severity error;5��    *   ?                  �                     �    *   B                 �                    5�_�   �   �           �   +   K    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f�C     �   *   ,   >      [        assert stimulus = "000001" report "Did not proceed to 1, count is " severity error;5��    *   K                  �                     �    *   M                 �                    �    *   O                  �                     �    *   N                 �                    �    *   P                                        �    *   O                  �                     �    *   N                 �                    �    *   N                 �                    �    *   N                 �                    5�_�   �   �           �   +   V    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f�Y     �   *   ,   >      l        assert stimulus = "000001" report "Did not proceed to 1, count is " & stimulus'image severity error;5��    *   V                                       5�_�   �   �           �   +   V    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f�Y     �   *   ,   >      k        assert stimulus = "000001" report "Did not proceed to 1, count is " & stimulusimage severity error;5��    *   V                                       5�_�   �   �           �   +   V    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f�[     �   *   ,   >      e        assert stimulus = "000001" report "Did not proceed to 1, count is " & stimulusseverity error;5��    *   V                                       5�_�   �   �           �   +   N    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f�p     �   *   ,   >      f        assert stimulus = "000001" report "Did not proceed to 1, count is " & stimulus severity error;5��    *   N                  �                     5�_�   �   �           �   +   Y    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f�u     �   *   ,   >      q        assert stimulus = "000001" report "Did not proceed to 1, count is " & to_integer(stimulus severity error;5��    *                     �      r       s       5�_�   �   �           �   +   X    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f�{     �   *   ,   >      r        assert stimulus = "000001" report "Did not proceed to 1, count is " & to_integer(stimulus) severity error;5��    *   X                                       5�_�   �   �           �   +   X    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f��     �   *   ,   >      x        assert stimulus = "000001" report "Did not proceed to 1, count is " & to_integersigned(stimulus) severity error;5��    *   X                                       5�_�   �   �           �   +   Y    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f��     �   *   ,   >      y        assert stimulus = "000001" report "Did not proceed to 1, count is " & to_integer(signed(stimulus) severity error;5��    *                     �      z       {       5�_�   �   �           �   +   j    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f��     �   *   ,   >      z        assert stimulus = "000001" report "Did not proceed to 1, count is " & to_integer(signed(stimulus)) severity error;5��    *   j                                       5�_�   �   �           �   +   l    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f��     �   *   ,   >      |        assert stimulus = "000001" report "Did not proceed to 1, count is " & to_integer(signed(stimulus))'' severity error;5��    *   k                                     5�_�   �   �           �   +   j    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f��     �   *   ,   >      �        assert stimulus = "000001" report "Did not proceed to 1, count is " & to_integer(signed(stimulus))'image severity error;5��    *   j                                       5�_�   �   �           �   +   j    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f��     �   *   ,   >              assert stimulus = "000001" report "Did not proceed to 1, count is " & to_integer(signed(stimulus))image severity error;5��    *   j                                       5�_�   �   �           �   +   j    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f��     �   *   ,   >      y        assert stimulus = "000001" report "Did not proceed to 1, count is " & to_integer(signed(stimulus))severity error;5��    *   j                                       5�_�   �   �   �       �   +   N    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f��     �   *   ,   >      z        assert stimulus = "000001" report "Did not proceed to 1, count is " & to_integer(signed(stimulus)) severity error;5��    *   N                  �                     5�_�   �   �           �   +   \    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f��     �   *   ,   >      �        assert stimulus = "000001" report "Did not proceed to 1, count is " & integer'image(to_integer(signed(stimulus)) severity error;5��    *                     �      �       �       5�_�   �   �           �   -   @    ����                                                                                                                                                                                                                                                                                                                            +   L       +   y       v   y    f��     �   ,   .   >      P        assert stimulus = "000010" report "Did not proceed to 2" severity error;�   -   .   >    5��    ,   A               .   �              .       5�_�   �   �           �   /   @    ����                                                                                                                                                                                                                                                                                                                            +   L       +   y       v   y    f�     �   .   0   >      P        assert stimulus = "000011" report "Did not proceed to 3" severity error;�   /   0   >    5��    .   A               .   8              .       5�_�   �   �           �   1   @    ����                                                                                                                                                                                                                                                                                                                            +   L       +   y       v   y    f�    �   0   2   >      P        assert stimulus = "000100" report "Did not proceed to 4" severity error;�   1   2   >    5��    0   A               .   �              .       5�_�   �   �           �   +   g    ����                                                                                                                                                                                                                                                                                                                            +   L       +   y       v   y    f�C     �   *   ,   >      �        assert stimulus = "000001" report "Did not proceed to 1, count is " & integer'image(to_integer(signed(stimulus))) severity error;5��    *   g                                     �    *   l                                     5�_�   �   �           �   -   \    ����                                                                                                                                                                                                                                                                                                                            +   L       +   y       v   y    f�R     �   ,   .   >      ~        assert stimulus = "000010" report "Did not proceed to 2" & integer'image(to_integer(signed(stimulus))) severity error;5��    ,   \                  �                     5�_�   �   �           �   /   \    ����                                                                                                                                                                                                                                                                                                                            +   L       +   y       v   y    f�Z     �   .   0   >      ~        assert stimulus = "000011" report "Did not proceed to 3" & integer'image(to_integer(signed(stimulus))) severity error;5��    .   \                  W                     5�_�   �   �           �   1   \    ����                                                                                                                                                                                                                                                                                                                            +   L       +   y       v   y    f�]   
 �   0   2   >      ~        assert stimulus = "000100" report "Did not proceed to 4" & integer'image(to_integer(signed(stimulus))) severity error;5��    0   \                  �                     5�_�   �   �   �       �   $        ����                                                                                                                                                                                                                                                                                                                            +   p       +   p       V   p    f��     �   #   %   ?              �   #   %   >    5��    #                      �              	       �    #                     �                     �    #   
                  �                     �    #   	                  �                     �    #                    �                    �    #                    �                    �    #                    �                    �    #                 2   �             2       5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            $          $          v       f�     �   #   %   ?      :        assert neg_condition report message severity note;5��    #                    �                    5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            $   "       $          v       f�     �   #   %   ?      2        assert false report message severity note;5��    #                     �                     5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            $   "       $          v       f�     �   #   %   ?      +        assert false report  severity note;5��    #                     �                     5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            $   "       $          v       f�     �   #   %   ?      -        assert false report "" severity note;5��    #                  	   �              	       5�_�   �   �           �   $   '    ����                                                                                                                                                                                                                                                                                                                            $   "       $          v       f�     �   #   %   ?      6        assert false report "batata e " severity note;5��    #   '                  �                     �    #   (                 �                    5�_�   �   �           �   $   *    ����                                                                                                                                                                                                                                                                                                                            $   "       $          v       f�     �   #   %   ?      9        assert false report "batata e " &  severity note;5��    #   *                  �                     5�_�   �   �           �   $   +    ����                                                                                                                                                                                                                                                                                                                            $   "       $          v       f�    �   #   %   ?      ;        assert false report "batata e " & "" severity note;5��    #   +                  �                     5�_�   �   �           �   .   >    ����                                                                                                                                                                                                                                                                                                                            ,   ?       ,   I       v   I    f��     �   -   /   ?      �        assert stimulus = "000010" report "Did not proceed to 2" & integer'image(to_integer(unsigned(stimulus))) severity error;�   .   /   ?    5��    -   ?                  �                     5�_�   �   �           �   0   >    ����                                                                                                                                                                                                                                                                                                                            0   H       0   H       v   H    f��     �   /   1   ?      �        assert stimulus = "000011" report "Did not proceed to 3" & integer'image(to_integer(unsigned(stimulus))) severity error;�   0   1   ?    5��    /   ?                  �                     5�_�   �   �           �   2   >    ����                                                                                                                                                                                                                                                                                                                            0   H       0   H       v   H    f��    �   1   3   ?      �        assert stimulus = "000100" report "Did not proceed to 4" & integer'image(to_integer(unsigned(stimulus))) severity error;�   2   3   ?    5��    1   ?                  1                     5�_�   �   �           �      	    ����                                                                                                                                                                                                                                                                                                                            0   H       0   H       v   H    f�B    �         ?      use IEEE.NUMERIC_STD.ALL;5��       	                 4                     �                         6                      �       
                  5                      �       	                 4                     �                         >                      �                         =                      �                         <                      �                         ;                      �                         :                      �                         9                      �                         8                      �                         7                      �                         6                      �       
                  5                      �       	                 4                     �       	                 4                     �       	                 4                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            0   H       0   H       v   H    f�M    �                use IEEE.STD_LOGIC_1164.ALL;5��                                                5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                            /   H       /   H       v   H    f�[    �   "   #          @        assert false report "batata e " & "arroz" severity note;5��    "                      �      A               5�_�   �   �           �   *   N    ����                                                                                                                                                                                                                                                                                                                            .   H       .   H       v   H    f�s     �   )   ,   =      �        assert stimulus = "000001" report "Did not proceed to 1, count is " & integer'image(to_integer(unsigned(stimulus))) severity error;5��    )   N                 �              	       5�_�   �   �           �   +   6    ����                                                                                                                                                                                                                                                                                                                            /   H       /   H       v   H    f�w     �   *   -   >      E        integer'image(to_integer(unsigned(stimulus))) severity error;5��    *   6                               	       5�_�   �   �           �   +   6    ����                                                                                                                                                                                                                                                                                                                            0   H       0   H       v   H    f�     �   *   -   ?      6        integer'image(to_integer(unsigned(stimulus))) 5��    *   6                                       �    *   :                               	       5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                            1   H       1   H       v   H    f��     �   +   -   @              5��    +                     %                     5�_�   �   �           �   ,   	    ����                                                                                                                                                                                                                                                                                                                            1   H       1   H       v   H    f��     �   +   -   @      
        ""5��    +   	               	   &              	       5�_�   �   �           �   *   *    ����                                                                                                                                                                                                                                                                                                                            1   H       1   H       v   H    f��     �   )   ,   @      N        assert stimulus = "000001" report "Did not proceed to 1, count is " & 5��    )   *                 �              	       5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                            2   H       2   H       v   H    f��     �   *   ,   A      ,        "Did not proceed to 1, count is " &    2integer'image(to_integer(unsigned(stimulus))) &LF&�   +   -   A      :        integer'image(to_integer(unsigned(stimulus))) &LF&5��    +                     �                     �    +                     �                     �    +                     �                     �    +                     �                     �    +                     �                     �    +                     �                     �    +                     �                     �    +                      �                     �    *   ,                  �                     5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                            1   H       1   H       v   H    f��     �   +   -   @              "Clock is "5��    +                     0                     5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                            +   ,       +   X       v   X    f��     �   +   -   @              "Clock is " �   ,   -   @    5��    +                  -   1              -       5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                            +   ,       +   X       v   X    f��     �   +   -   @      A        "Clock is " integer'image(to_integer(unsigned(stimulus)))5��    +                     0                     5�_�   �   �           �   ,   8    ����                                                                                                                                                                                                                                                                                                                            +   ,       +   X       v   X    f��    �   +   -   @      C        "Clock is " & integer'image(to_integer(unsigned(stimulus)))5��    +   8                 U                    5�_�   �   �           �   /   *    ����                                                                                                                                                                                                                                                                                                                            /   *       /   {       v   {    f��     �   .   1   @      �        assert stimulus = "000010" report "Did not proceed to 2, count is " & integer'image(to_integer(unsigned(stimulus))) severity error;5��    .   *       R           �      R               �    .   *                 �              	       5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            ,          +          V       f��     �   /   2   A    �   /   0   A    5��    /                      �              �       5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                            ,          +          V       f��     �   -   /   C    5��    -                      t              	       �    -                     {                     �    -                     z                     �    -                     y                     �    -                     x                     �    -                     w                     �    -                     v                     �    -                     u                     �    -                      t                     5�_�   �   �           �   4        ����                                                                                                                                                                                                                                                                                                                            ,          +          V       f��     �   3   5   D    5��    3                      u              	       �    3                     |                     �    3                     {                     �    3                     z                     �    3                     y                     �    3                     x                     �    3                     w                     �    3                     v                     �    3                      u                     5�_�   �   �           �   7        ����                                                                                                                                                                                                                                                                                                                            ,          +          V       f��     �   6   8   E    5��    6                      !              	       �    6                     (                     �    6                     '                     �    6                     &                     �    6                     %                     �    6                     $                     �    6                     #                     �    6                     "                     �    6                      !                     5�_�   �   �   �       �   :        ����                                                                                                                                                                                                                                                                                                                            ,          +          V       f��     �   9   ;   F    5��    9                      �              	       �    9                     �                     �    9                     �                     �    9                     �                     �    9                     �                     �    9                     �                     �    9                     �                     �    9                     �                     �    9                      �                     5�_�   �   �           �   6   *    ����                                                                                                                                                                                                                                                                                                                            6   *       6   {       v   {    f��     �   5   8   G      �        assert stimulus = "000011" report "Did not proceed to 3, count is " & integer'image(to_integer(unsigned(stimulus))) severity error;5��    5   *       R           �      R               �    5   *                 �              	       5�_�   �   �           �   6       ����                                                                                                                                                                                                                                                                                                                            2          1          V       f�     �   6   9   H    �   6   7   H    5��    6                      �              �       5�_�   �   �           �   1       ����                                                                                                                                                                                                                                                                                                                            2          1          V       f�     �   0   2   J      ^        "Did not proceed to 1, count is " & integer'image(to_integer(unsigned(stimulus))) &LF&5��    0                    �                    5�_�   �   �           �   7       ����                                                                                                                                                                                                                                                                                                                            2          1          V       f�	     �   6   8   J      ^        "Did not proceed to 1, count is " & integer'image(to_integer(unsigned(stimulus))) &LF&5��    6                    �                    5�_�   �   �           �   <   *    ����                                                                                                                                                                                                                                                                                                                            <   *       <   {       v   {    f�     �   ;   >   J      �        assert stimulus = "000100" report "Did not proceed to 4, count is " & integer'image(to_integer(unsigned(stimulus))) severity error;5��    ;   *       R           �      R               �    ;   *                 �              	       5�_�   �   �           �   <       ����                                                                                                                                                                                                                                                                                                                            8          7          V       f�     �   <   ?   K    �   <   =   K    5��    <                      �              �       5�_�   �   �           �   =       ����                                                                                                                                                                                                                                                                                                                            8          7          V       f�!    �   <   >   M      ^        "Did not proceed to 3, count is " & integer'image(to_integer(unsigned(stimulus))) &LF&5��    <                    �                    5�_�   �   �           �   >       ����                                                                                                                                                                                                                                                                                                                            8          7          V       f�4     �   =   ?   M      >        "Clock is " & integer'image(to_integer(unsigned(clk)))5��    =                    6                    5�_�   �   �           �   >        ����                                                                                                                                                                                                                                                                                                                            8          7          V       f�9    �   =   ?   M      :        "Clock is " & bit'image(to_integer(unsigned(clk)))5��    =                     @                    5�_�   �   �           �   8   "    ����                                                                                                                                                                                                                                                                                                                            8          7          V       f�?     �   8   :   M    �   8   9   M    5��    8                      ^              %       5�_�   �   �   �       �   2       ����                                                                                                                                                                                                                                                                                                                            8          7          V       f�A     �   2   4   N    �   2   3   N    5��    2                      ]              %       5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                            9          8          V       f�C     �   ,   .   O    �   -   .   O    5��    ,                      \              %       5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                            :          9          V       f�D     �   +   ,          >        "Clock is " & integer'image(to_integer(unsigned(clk)))5��    +                            ?               5�_�   �   �           �   2       ����                                                                                                                                                                                                                                                                                                                            9          8          V       f�F     �   1   2          >        "Clock is " & integer'image(to_integer(unsigned(clk)))5��    1                            ?               5�_�   �   �           �   8       ����                                                                                                                                                                                                                                                                                                                            8          7          V       f�G    �   7   8          >        "Clock is " & integer'image(to_integer(unsigned(clk)))5��    7                      �      ?               5�_�   �   �   �       �      -    ����                                                                                                                                                                                                                                                                                                                            8          7          V       f�     �         M      L    signal stimulus : bit_vector(5 downto 0) := "000000";  -- Input stimulus5��       -                  i                     �       ,                  h                     5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            8          7          V       f�    �   &   '                   -- stimulus <= "000000";5��    &                      F      !               5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            7          6          V       f
     �         L      /    signal reset : bit := '0';  -- Reset signal5��                        '                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            7          6          V       f     �         L      /    signal reset : bit := '1';  -- Reset signal5��                                            5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            7          6          V       f     �         L      @    signal stimulus : bit_vector(5 downto 0);  -- Input stimulus5��                        E                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            7          6          V       f     �         L                  rst => reset,5��                                            5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            7          6          V       f     �         L                  count => stimulus5��                        0                    �                         4                     �                        3                    5�_�   �   �           �   )       ����                                                                                                                                                                                                                                                                                                                            7          6          V       f     �   (   *   L      *        assert stimulus = "000001" report 5��    (                    k                    5�_�   �   �           �   *        ����                                                                                                                                                                                                                                                                                                                            *          ?           V       f+     �   ;   =          ^        "Did not proceed to 4, count is " & integer'image(to_integer(unsigned(stimulus))) &LF&�   :   <          *        assert stimulus = "000100" report �   5   7          ^        "Did not proceed to 3, count is " & integer'image(to_integer(unsigned(stimulus))) &LF&�   4   6          *        assert stimulus = "000011" report �   /   1          ^        "Did not proceed to 2, count is " & integer'image(to_integer(unsigned(stimulus))) &LF&�   .   0          *        assert stimulus = "000010" report �   )   +   L      ^        "Did not proceed to 1, count is " & integer'image(to_integer(unsigned(stimulus))) &LF&5��    )   N                 �                    �    .                    L                    �    /   N                 �                    �    4                    -                    �    5   N                 �                    �    :                                        �    ;   N                 u                    5�_�   �   �           �   B       ����                                                                                                                                                                                                                                                                                                                            *          ?           V       fJ     �   A   B                   -- stimulus <= "001011";5��    A                      �      !               5�_�   �   �           �   G       ����                                                                                                                                                                                                                                                                                                                            B          G          V       fN     �   A   H   K      )        -- reset <= '1';  -- Assert reset   :        -- wait for CLOCK_PERIOD;  -- Hold reset for 20 ns   L        -- assert stimulus = "000000" report "Did not reset" severity error;   +        -- reset <= '0';  -- Deassert reset   :        -- wait for CLOCK_PERIOD;  -- Hold reset for 20 ns   N        -- assert stimulus = "000001" report "Did not proceed" severity error;5��    A                     �      h      V      5�_�   �   �           �   B       ����                                                                                                                                                                                                                                                                                                                            B          G          V       fR     �   A   C   K      &        reset <= '1';  -- Assert reset5��    A                    �                    5�_�   �   �           �   E       ����                                                                                                                                                                                                                                                                                                                            B          G          V       fT     �   D   F   K      (        reset <= '0';  -- Deassert reset5��    D                    �                    �    D   	                 �                    5�_�   �   �           �   D       ����                                                                                                                                                                                                                                                                                                                            B          G          V       fX     �   C   E   K      I        assert stimulus = "000000" report "Did not reset" severity error;5��    C                    M                    5�_�   �   �           �   G       ����                                                                                                                                                                                                                                                                                                                            B          G          V       f[    �   F   H   K      K        assert stimulus = "000001" report "Did not proceed" severity error;5��    F                    �                    5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                            B          G          V       f     �   %   '   K              wait for CLOCK_PERIOD;5��    %                     :                     5�_�   �   �           �   &        ����                                                                                                                                                                                                                                                                                                                            B          G          V       f�     �   &   (   L              �   &   (   K    5��    &                      @              	       �    &                     H                     �    &   	                  I                     �    &                    H                    �    &                    H                    �    &                    H                    �    &                 2   H             2       5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            '          '          v       f�     �   &   (   L      :        assert neg_condition report message severity note;5��    &                    O                    5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            '   "       '          v       f�     �   &   )   L      2        assert false report message severity note;5��    &                    \                    �    &                     ]                     �    &                     \                     �    &                     [                     �    &                   [             	       5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                            '   "       '          v       f�     �   ,   -          $        "Clock is " & bit'image(clk)5��    ,                            %               5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                            '   "       '          v       f�     �   '   )   L    �   (   )   L    5��    '                      \              %       5�_�   �   �           �   -   V    ����                                                                                                                                                                                                                                                                                                                            '   "       '          v       f�     �   ,   .   M      [        "Did not proceed to 1, count is " & integer'image(to_integer(unsigned(count))) &LF&5��    ,   V                  6                     5�_�   �   �           �   2   V    ����                                                                                                                                                                                                                                                                                                                            '   "       '          v       f�     �   1   3   M      [        "Did not proceed to 2, count is " & integer'image(to_integer(unsigned(count))) &LF&5��    1   V                  �                     5�_�   �   �           �   3   #    ����                                                                                                                                                                                                                                                                                                                            '   "       '          v       f�     �   2   3          $        "Clock is " & bit'image(clk)5��    2                      �      %               5�_�   �   �           �   7   W    ����                                                                                                                                                                                                                                                                                                                            '   "       '          v       f�     �   6   8   L      [        "Did not proceed to 3, count is " & integer'image(to_integer(unsigned(count))) &LF&5��    6   W                  �                     5�_�   �   �           �   7   V    ����                                                                                                                                                                                                                                                                                                                            '   "       '          v       f�     �   6   8   L      W        "Did not proceed to 3, count is " & integer'image(to_integer(unsigned(count))) 5��    6   V                  �                     5�_�   �   �           �   8   #    ����                                                                                                                                                                                                                                                                                                                            '   "       '          v       f�     �   7   8          $        "Clock is " & bit'image(clk)5��    7                      �      %               5�_�   �   �           �   <   W    ����                                                                                                                                                                                                                                                                                                                            '   "       '          v       f�     �   ;   =   K      [        "Did not proceed to 4, count is " & integer'image(to_integer(unsigned(count))) &LF&5��    ;   W                  \                     5�_�   �   �           �   =   #    ����                                                                                                                                                                                                                                                                                                                            '   "       '          v       f�    �   <   =          $        "Clock is " & bit'image(clk)5��    <                      ]      %               5�_�   �   �           �   )        ����                                                                                                                                                                                                                                                                                                                            &          )          V       f�     �   )   .   J    �   )   *   J    5��    )                      �              {       5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                            &          )          V       f�    �   -   2   N    �   -   .   N    5��    -                                    {       5�_�   �   �   �       �          ����                                                                                                                                                                                                                                                                                                                            &          )          V       f	�     �         S          �         R    5��                          �                     �                         �                     �                         �                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            '          *          V       f	�     �         S          rst <= 5��                         �                     5�_�   �              �          ����                                                                                                                                                                                                                                                                                                                            '          *          V       f	�     �         S          rst <= ''5��                         �                     5�_�   �                       ����                                                                                                                                                                                                                                                                                                                            '          *          V       f	�     �         S          rst <= '1'5��                         �                     �                         �                     5�_�                         ����                                                                                                                                                                                                                                                                                                                            '          *          V       f	�     �         S          rst <= '1', 5��                         �                     5�_�                        ����                                                                                                                                                                                                                                                                                                                            '          *          V       f	�     �         S          rst <= '1', ''5��                         �                     5�_�                        ����                                                                                                                                                                                                                                                                                                                            '          *          V       f	�     �         S          rst <= '1', '0'5��                         �                     �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    �                         �                     5�_�                        ����                                                                                                                                                                                                                                                                                                                            '          *          V       f	�     �         S          rst <= '1', '0' after5��                         �                     5�_�                        ����                                                                                                                                                                                                                                                                                                                            '          *          V       f	�     �         S          rst <= '1', '0' after()5��                         �                     �                        �                    �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    5�_�                    &    ����                                                                                                                                                                                                                                                                                                                            '          *          V       f	�     �         S      &    rst <= '1', '0' after CLOCK_PERIOD5��       &                  �                     5�_�                 $        ����                                                                                                                                                                                                                                                                                                                            $   &       &   &       V   &    f	�     �   #   $          +        -- Apply stimulus to the DUT inputs   6        -- You can control the timing of stimulus here   C        -- For example, change the stimulus value every clock cycle5��    #                      �      �               5�_�    	             $   !    ����                                                                                                                                                                                                                                                                                                                            $   &       $   &       V   &    f	�     �   #   %   Q              �   #   %   P    5��    #                      �              	       �    #                     �                     �    #                     �                     �    #                     �                     �    #                     �                     �    #                     �                     �    #                     �                     �    #                    �                    �    #                 
   �             
       5�_�    
          	   $       ����                                                                                                                                                                                                                                                                                                                            %   &       %   &       V   &    f	�     �   #   %   Q              wait until rst = 5��    #                     �                     5�_�  	            
   $       ����                                                                                                                                                                                                                                                                                                                            %   &       %   &       V   &    f	�     �   #   %   Q              wait until rst = ''5��    #                     �                     5�_�  
               $       ����                                                                                                                                                                                                                                                                                                                            %   &       %   &       V   &    f	�     �   #   %   Q              wait until rst = '0'5��    #                     �                     5�_�                 $       ����                                                                                                                                                                                                                                                                                                                            %   &       %   &       V   &    f	�    �   $   &   Q    5��    $                      �              	       �    $                     �                     �    $                     �                     �    $                     �                     �    $                     �                     �    $                     �                     �    $                     �                     �    $                     �                     �    $                      �                     5�_�                       ����                                                                                                                                                                                                                                                                                                                            &           2           V        f    �                '    rst <= '1', '0' after CLOCK_PERIOD;5��                          �      (               5�_�                 #        ����                                                                                                                                                                                                                                                                                                                            %           %           V        f+    �   "   #                  wait until rst = '0';5��    "                      v                     5�_�                        ����                                                                                                                                                                                                                                                                                                                                       P           V        f�    �         P      -    signal rst : bit := '1';  -- Reset signal5��                        %                    5�_�                      ����                                                                                                                                                                                                                                                                                                                                       P           V        f     �         Q          �         Q    �         P    5��                          �                     �                  	      �              �       5�_�                         ����                                                                                                                                                                                                                                                                                                                                                          fL     �         Z      clk_process: process5��                          �                     5�_�                       ����                                                                                                                                                                                                                                                                                                                                                          fP     �         Z      begin5��                                               5�_�                        ����                                                                                                                                                                                                                                                                                                                                                       fT     �         Z          wait for CLOCK_PERIOD / 2;       while true loop           clk <= not clk;   "        wait for CLOCK_PERIOD / 2;       end loop;�         Z          clk <= '0';5��                                              �                         -                     �                         P                     �                         h                     �                         �                     �                         �                     5�_�                         ����                                                                                                                                                                                                                                                                                                                                                       fW     �         Z      end process clk_process;5��                          �                     5�_�                         ����                                                                                                                                                                                                                                                                                                                                                V       f`     �             
       -- Clock process       clk_process: process   	    begin           clk <= '0';   "        wait for CLOCK_PERIOD / 2;           while true loop               clk <= not clk;   &            wait for CLOCK_PERIOD / 2;           end loop;       end process clk_process;5��           
               �      �               5�_�                         ����                                                                                                                                                                                                                                                                                                                                                V       fb     �      !   P    �         P    5��                   
       �              �       5�_�                        ����                                                                                                                                                                                                                                                                                                                                                V       fe    �                (    clk <= clk after (CLOCK_PERIOD / 2);5��                                )               5�_�                 -        ����                                                                                                                                                                                                                                                                                                                                                V       fu    �   ,   -          "        wait for CLOCK_PERIOD / 2;           assert false report   $        "Clock is " & bit'image(clk)           severity note;   "        wait for CLOCK_PERIOD / 2;           assert false report   $        "Clock is " & bit'image(clk)           severity note;   "        wait for CLOCK_PERIOD / 2;           assert false report   $        "Clock is " & bit'image(clk)           severity note;    5��    ,                      G      r              5�_�               I        ����                                                                                                                                                                                                                                                                                                                                                V       f�     �   I   K   L    �   I   J   L    5��    I                      �              =       5�_�                  J       ����                                                                                                                                                                                                                                                                                                                                                V       f�     �   J   L   M    5��    J                      �              	       �    J                      �                     5�_�    !              J   !    ����                                                                                                                                                                                                                                                                                                                                                V       f�     �   I   K   N      <        assert false report "EOT ch function" severity note;5��    I   !                  �                     5�_�     "          !   J   !    ����                                                                                                                                                                                                                                                                                                                                                V       f�     �   I   K   N      :        assert false report "EOT  function" severity note;5��    I   !                  �                     5�_�  !  $          "   J   !    ����                                                                                                                                                                                                                                                                                                                                                V       f�     �   I   K   N      9        assert false report "EOT function" severity note;5��    I   !                 �                    5�_�  "  %  #      $   +       ����                                                                                                                                                                                                                                                                                                                                                V       f�     �   +   -   N    5��    +                      F                     �    +                     F                    �    +                     G                     �    +                      F                     5�_�  $  &          %   ,        ����                                                                                                                                                                                                                                                                                                                                                V       f�     �   ,   .   O    �   ,   -   O    5��    ,                      G              7       5�_�  %  '          &   -       ����                                                                                                                                                                                                                                                                                                                                                V       f�    �   ,   .   P      6        assert false report "EOT count" severity note;5��    ,                    d                    5�_�  &  (          '          ����                                                                                                                                                                                                                                                                                                                                                  V        f�8     �   
      P      U            count : out bit_vector(5 downto 0)       -- 6-bit count output (64 steps)5��    
                    5                    5�_�  '  )          (   0       ����                                                                                                                                                                                                                                                                                                                            0          0          v       f�E     �   /   1   P      '        assert count = "000001" report 5��    /                    �                    5�_�  (  *          )          ����                                                                                                                                                                                                                                                                                                                            0          0          v       f�R     �         P      =    signal count : bit_vector(5 downto 0);  -- Input stimulus5��                        >                    5�_�  )  +          *   5       ����                                                                                                                                                                                                                                                                                                                            0          0          v       f�[     �   4   6   P      '        assert count = "000010" report 5��    4          	          G      	              5�_�  *  ,          +   :       ����                                                                                                                                                                                                                                                                                                                            0          0          v       f�b     �   9   ;   P      '        assert count = "000011" report 5��    9          	          �      	              5�_�  +  -          ,   ?       ����                                                                                                                                                                                                                                                                                                                            0          0          v       f�f     �   >   @   P      '        assert count = "000100" report 5��    >          	          �      	              5�_�  ,  .          -   G       ����                                                                                                                                                                                                                                                                                                                            0          0          v       f�j     �   F   H   P      F        assert count = "000000" report "Did not reset" severity error;5��    F          	          �      	              5�_�  -              .   J       ����                                                                                                                                                                                                                                                                                                                            0          0          v       f�n     �   I   K   P      H        assert count = "000001" report "Did not proceed" severity error;5��    I          	          U      	              5�_�  "          $  #   +       ����                                                                                                                                                                                                                                                                                                                                                V       f�     �   +   ,   N    �   +   ,   N      6        assert false report "EOT count" severity note;5��    +                      F              7       5�_�               L       ����                                                                                                                                                                                                                                                                                                                                                V       fE     �   K   L   L          �   K   M   M      end dut;5��    K                      �                     �    K                      �                     �    K                      �                     �    K                     �                     5�_�                 L       ����                                                                                                                                                                                                                                                                                                                                                V       f/     �   L   M           �   L   N          end dut;5��    L                      �                     �    L                      �                     5�_�                        ����                                                                                                                                                                                                                                                                                                                                                          fN     �         Z      beg  in5��                                              5�_�                        ����                                                                                                                                                                                                                                                                                                                                       Q           V        f     �         P       5��                          �                     �                         �                     �                         �                     �                         �                     �                          �                     5�_�                 &        ����                                                                                                                                                                                                                                                                                                                            &           &           V        f	�     �   %   4        5��    %                      �      �              5�_�   �   �   �   �   �      	    ����                                                                                                                                                                                                                                                                                                                            '          *          V       f	|     �         R          �         S    �         S      !    reset <= '1', '0' after 5 ns;5��                          :                     �                         >                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            '          *          V       f	�     �         S      &    signal rst <= '1', '0' after 5 ns;5��                     
   >             
       5�_�   �   �   �       �          ����                                                                                                                                                                                                                                                                                                                            '          *          V       f	�     �         S      ,    signal rst : bit := '1', '0' after 5 ns;5��                        I                    5�_�   �               �          ����                                                                                                                                                                                                                                                                                                                            '          *          V       f	�     �         S      ,    signal rst : bit := '1'; '0' after 5 ns;5��                        U                    5�_�   �           �   �          ����                                                                                                                                                                                                                                                                                                                            &          )          V       f	�     �              5��                                .               5�_�   �   �       �   �      	    ����                                                                                                                                                                                                                                                                                                                            &          )          V       f	"     �         R          dut: work.counter_6bit5��       	                  �                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            &          )          V       f	$     �         R          dut: work.counter_6bit()5��                         �                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            &          )          V       f	-     �         R          dut: work.counter_6bit(rtl)5��                         �                     5�_�   �               �      	    ����                                                                                                                                                                                                                                                                                                                            &          )          V       f	7     �         R      &    dut: entity work.counter_6bit(rtl)5��       	                  �                     �                        �                    5�_�   �           �   �          ����                                                                                                                                                                                                                                                                                                                            7          6          V       f�     �              5��                          <      M               5�_�   �           �   �   9       ����                                                                                                                                                                                                                                                                                                                            8          7          V       f�?     �   9   :   N    �   9   :   N      $        "Clock is " & bit'image(clk)5��    9                      �              %       5�_�   �           �   �   :        ����                                                                                                                                                                                                                                                                                                                            ,          +          V       f��     �   :   ;   F       5��    :                      �              	       �    :                     �                     �    :                     �                     �    :                     �                     �    :                     �                     �    :                     �                     �    :                     �                     �    :                     �                     �    :                      �                     5�_�   �       �   �   �   +   p    ����                                                                                                                                                                                                                                                                                                                            +   L       +   y       v   y    f��   	 �   *   ,   >      �        assert stimulus = "000001" report "Did not proceed to 1, count is " & integer'image(to_integer(unsigned(count))) severity error;5��    *   p                                      �    *   q                  !                     �    *   p                                      �    *   s                  #                     �    *   r                  "                     �    *   q                  !                     �    *   p                                      �    *   t                  $                     �    *   s                  #                     �    *   r                  "                     �    *   q                  !                     �    *   p                                      �    *   p                                      �    *   p                                      5�_�   �           �   �   +   g    ����                                                                                                                                                                                                                                                                                                                            +   L       +   y       v   y    f�t     �   *   ,   >      �        assert stimulus = "000001" report "Did not proceed to 1, count is " & integer'image(to_integer(to_unsigned(stimulus))) severity error;5��    *   g                                       5�_�   �           �   �   +   Y    ����                                                                                                                                                                                                                                                                                                                            4           :           V        f��     �   *   ,   >      }        assert stimulus = "000001" report "Did not proceed to 1, count is " & to_integer(to_signed(stimulus)) severity error;5��    *   Y                  	                     5�_�   q   s       v   r          ����                                                                                                                                                                                                                                                                                                                            8          8           v        f��     �              5��                                                5�_�   r   t           s          ����                                                                                                                                                                                                                                                                                                                            7          7           v        f��     �              5��                                                5�_�   s   u           t           ����                                                                                                                                                                                                                                                                                                                            6          6           v        f��     �               5��                                                  5�_�   t               u           ����                                                                                                                                                                                                                                                                                                                            5          5           v        f��     �               5��                                                  5�_�   =           ?   >   C       ����                                                                                                                                                                                                                                                                                                                            5          4          V       f�      �   B   D   G       5��    B           (           g      (               5�_�   &           (   '   0       ����                                                                                                                                                                                                                                                                                                                            
                           f�D     �   /   0   C       5��    /                      z              	       �    /                      z                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                         +       v   (    f�     �         =       5��                          a                      �                          a                      �                          a                      5�_�              	             ����                                                                                                                                                                                                                                                                                                                                                V       f ǵ     �         =      entity counert is end;5��                         Q                      5�_�                          ����                                                                                                                                                                                                                                                                                                                                                V       f Ǭ     �              �         ;       5��                          j       4               �               #           F       #               5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f Ǧ     �         =      architecture Behavioral of  is5��                         �                      5��