Vim�UnDo� 
v��3����3��[�SPK�9�;��!6.�P�=   W                                   f(>.    _�                             ����                                                                                                                                                                                                                                                                                                                                                             f(=�     �                   �               5��                                         =      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f(=�    �                  5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f(>,     �               5��                          =                     5�_�                             ����                                                                                                                                                                                                                                                                                                                                                             f(>-    �               �               5��                   :       >              �      5��