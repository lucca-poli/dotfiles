Vim�UnDo� An���p�0M�q��^�/�JA��A��-�T�   �   .                                state <= idle;   �          n       n   n   n    f(��   	 _�                     v       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   u   w        		  shift: out bit;5��    u                     �	                     5�_�                    u   #    ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   t   v        #        done, parity_bit: out bit;5��    t   "                  �	                     5�_�                    v       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   u   w        		  shift: out bit;5��    u                     �	                     5�_�                    w       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   v   x        4		  internal_data: out bit_vector(WIDTH-1 downto 0);5��    v                     �	                     5�_�                    g       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   f   h            5��    f                      P                     5�_�                    f       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   e   g        	 new_clk <= clk_out;5��    e                     N                     5�_�                    e       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   d   f        	 5��    d                     7                     5�_�      	              d       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   c   e            end process timing;5��    c                     3                     5�_�      
           	   c       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   b   d                end if;5��    b                                          5�_�   	              
   b       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   a   c        				end if;5��    a                     	                     5�_�   
                 a       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   `   b        					CNT <= CNT + 1;5��    `                     �                     5�_�                    `   	    ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   _   a        					else5��    _                     �                     5�_�                    _       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   ^   `        					CLK_OUT <= not CLK_OUT;5��    ^                     �                     5�_�                    ^       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   ]   _        					CNT <= 0;5��    ]                     �                     5�_�                    ]       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   \   ^        				if cnt = MAX_CNT then5��    \                     �                     5�_�                    \   $    ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   [   ]        $        if rising_edge(clk_in) then5��    [   #                  �                     5�_�                    [   
    ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   Z   \        
    begin5��    Z   	                  n                     5�_�                    Z       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   Y   [            timing: process(clk_in)5��    Y                     c                     5�_�                    Y       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   X   Z            5��    X                     F                     5�_�                    X       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   W   Y        begin5��    W                     @                     5�_�                    W       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   V   X            5��    V                     9                     5�_�                    V   )    ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   U   W        )    constant MAX_CNT: natural := factor;5��    U   (                  3                     5�_�                    U       ����                                                                                                                                                                                                                                                                                                                                                             f(;�     �   T   V        	 signal CLK_OUT: bit := '0';5��    T                     	                     5�_�                    T       ����                                                                                                                                                                                                                                                                                                                                                             f(<      �   S   U            signal CNT: natural := 0;5��    S                     �                     5�_�                    S       ����                                                                                                                                                                                                                                                                                                                                                             f(<     �   R   T        5��    R                      �                     5�_�                    R        ����                                                                                                                                                                                                                                                                                                                                                             f(<    �   Q   S         architecture rtl of slow_clk is5��    Q                     �                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                      C          V       f(=G     �             &   library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity counter_generic is       generic(           MAX_COUNT: natural       );   
    port (   J        clk, rst, start: in bit;                            -- Clock input           done: out bit;   B        count : out natural       -- 6-bit count output (64 steps)       );   end counter_generic;       -architecture Behavioral of counter_generic is   !    signal counter: natural := 0;       begin          &    counting: process(clk, rst, start)   	    begin           if rst = '1' then               counter <= 0;               done <= '0';   #        elsif rising_edge(clk) then   )            if counter = MAX_COUNT-1 then                   done <= '1';                   counter <= 0;               end if;   \            if (counter > 0 and counter < MAX_COUNT-1) or (start = '1' and counter = 0) then   '                counter <= counter + 1;               end if;           end if;       end process counting;           count <= counter;          end architecture;5��           &               >      �              5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       f(=P     �          �      library IEEE;5��                         L                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       f(=Q     �      !   �      use IEEE.NUMERIC_BIT.all;5��                         f                     5�_�                    !       ����                                                                                                                                                                                                                                                                                                                                                V       f(=R     �       "   �      5��                           g                     5�_�                     "       ����                                                                                                                                                                                                                                                                                                                                                V       f(=S     �   !   #   �      entity slow_clk is5��    !                     z                     5�_�      !               #       ����                                                                                                                                                                                                                                                                                                                                                V       f(=T     �   "   $   �      	 generic(5��    "   
                  �                     5�_�       "           !   $       ����                                                                                                                                                                                                                                                                                                                                                V       f(=U     �   #   %   �      			factor: natural5��    #                     �                     5�_�   !   #           "   %       ����                                                                                                                                                                                                                                                                                                                                                V       f(=W     �   $   &   �       );5��    $                     �                     5�_�   "   $           #   #       ����                                                                                                                                                                                                                                                                                                                                                V       f(=Y     �   "   $   �      
	 generic(5��    "                     |                     5�_�   #   %           $   %       ����                                                                                                                                                                                                                                                                                                                                                V       f(=\     �   $   &   �       );5��    $                     �                     5�_�   $   &           %   &       ����                                                                                                                                                                                                                                                                                                                                                V       f(=]     �   %   '   �          port (5��    %   
                  �                     5�_�   %   '           &   '       ����                                                                                                                                                                                                                                                                                                                                                V       f(=^     �   &   (   �              clk_in: in bit;5��    &                     �                     5�_�   &   (           '   (       ����                                                                                                                                                                                                                                                                                                                                                V       f(=_     �   '   )   �              new_clk: out bit5��    '                     �                     5�_�   '   )           (   )       ����                                                                                                                                                                                                                                                                                                                                                V       f(=`     �   (   *   �          );5��    (                     �                     5�_�   (   *           )   *       ����                                                                                                                                                                                                                                                                                                                                                V       f(=f     �   )   +   �      end entity slow_clk;5��    )                     �                     5�_�   )   +           *   +       ����                                                                                                                                                                                                                                                                                                                                                V       f(=g     �   *   ,   �      5��    *                      �                     5�_�   *   ,           +           ����                                                                                                                                                                                                                                                                                                                                       B           V        f(=o     �             $   library IEEE;   use IEEE.NUMERIC_BIT.all;       entity slow_clk is   		generic(   			factor: natural       );   
    port (           clk_in: in bit;           new_clk: out bit       );   end entity slow_clk;       architecture rtl of slow_clk is           signal CNT: natural := 0;   	 signal CLK_OUT: bit := '0';   (    constant MAX_CNT: natural := factor;          begin              timing: process(clk_in)   	    begin   #        if rising_edge(clk_in) then   				if cnt = MAX_CNT then   					CNT <= 0;   					CLK_OUT <= not CLK_OUT;   				else   					CNT <= CNT + 1;   				end if;           end if;       end process timing;   	    	 new_clk <= clk_out;       end architecture rtl;5��           $               ?      a              5�_�   +   -           ,           ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �                 library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity shift_reg8 is   
    port (   !        rst, clk, enable: in bit;           data: in bit;   %        q: out bit_vector(7 downto 0)       );   end entity;       &architecture Behavior of shift_reg8 is   =   signal vector: bit_vector(7 downto 0) := (others => '0');        begin              process(rst, clk)   	    begin           if rst = '1' then   &            vector <= (others => '0');   4        elsif rising_edge(clk) and enable = '1' then   0            vector <= data & vector(7 downto 1);           end if;       end process;           q <= vector;          end architecture;5��                                   =              5�_�   ,   1           -           ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �                      5��                                                  5�_�   -   2   .       1   �       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   �   �   �      	 5��    �                     �                     5�_�   1   3           2   �       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   �   �   �          end process;5��    �                     �                     5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �                2		internal_data: out bit_vector(WIDTH-1 downto 0);5��                          @      3               5�_�   3   5           4   �       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   �   �          	 internal_data <= word;5��    �                      �                     5�_�   4   6           5   �       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   �   �          	 shift <= shift_data;5��    �                      �                     5�_�   5   7           6   �        ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   �   �          	 5��    �                      �                     5�_�   6   8           7          ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �                		shift: out bit;5��                          .                     5�_�   7   9           8   .       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   -   /   �              new_clk: out bit5��    -                     k                     5�_�   8   :           9   -       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   ,   .   �              clk_in: in bit;5��    ,                     Q                     5�_�   9   ;           :   ,       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   +   -   �          port (5��    +   
                  8                     5�_�   :   <           ;   +       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   *   ,   �      	 );5��    *                     ,                     5�_�   ;   =           <   *       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   )   +   �      			factor: natural5��    )                     &                     5�_�   <   >           =   )       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   (   *   �      			generic(5��    (                                          5�_�   =   ?           >   (       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   '   )   �          component slow_clk5��    '                                          5�_�   >   A           ?   )       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   (   *   �      			generic(5��    (                                          5�_�   ?   B   @       A   +       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   *   ,   �      	 );5��    *                     &                     5�_�   A   C           B   ,       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   +   -   �      
    port (5��    +                     0                     5�_�   B   D           C   -       ����                                                                                                                                                                                                                                                                                                                            -          .                 f(=�     �   -   /   �              new_clk: out bit�   ,   .   �              clk_in: in bit;5��    ,                     C                     �    -                     _                     5�_�   C   E           D   /       ����                                                                                                                                                                                                                                                                                                                            -          .                 f(=�     �   .   0   �          );5��    .                     x                     5�_�   D   F           E   �       ����                                                                                                                                                                                                                                                                                                                            -          .                 f(=�     �   �   �              5��    �                      �                     5�_�   E   H           F   �       ����                                                                                                                                                                                                                                                                                                                                                             f(=�    �   �   �   �    5��    �                      �                     �    �                      �                     �    �                      �                     5�_�   F   I   G       H   I       ����                                                                                                                                                                                                                                                                                                                                                             f(m]     �   H   J   �          clocking: slow_clk5��    H                                          5�_�   H   M           I   J       ����                                                                                                                                                                                                                                                                                                                                                             f(m_    �   I   K   �      			generic map(1)5��    I                                          5�_�   I   N   J       M          ����                                                                                                                                                                                                                                                                                                                            :           ;           V        f(�-     �         �      1        clock, reset, start, serial_data: in bit;5��                         �                      5�_�   M   O           N          ����                                                                                                                                                                                                                                                                                                                            :           ;           V        f(�K     �                        PARITY: natural := 1;           CLOCK_MUL: natural := 45��                          �       >               5�_�   N   P           O          ����                                                                                                                                                                                                                                                                                                                            8           9           V        f(�L     �                "        POLARITY: boolean := TRUE;5��                          J       #               5�_�   O   Q           P          ����                                                                                                                                                                                                                                                                                                                            7           8           V        f(�L     �         �              WIDTH: natural := 7;5��                         e                      5�_�   P   R           Q   d       ����                                                                                                                                                                                                                                                                                                                            7           8           V        f(�R     �   c   e   �      A                        if start = '1' and serial_data = '0' then5��    c                     
                     5�_�   Q   S           R   �       ����                                                                                                                                                                                                                                                                                                                            7           8           V        f(�W    �   �   �   �      E                            if start = '1' and serial_data = '0' then5��    �                     G                     5�_�   R   T           S          ����                                                                                                                                                                                                                                                                                                                                                V       f(��     �         �      entity serial_in is5��              	          0       	              5�_�   S   [           T          ����                                                                                                                                                                                                                                                                                                                                                V       f(��    �         �      'architecture Behavioral of serial_in is5��              	          +      	              �                         0                    5�_�   T   \   X       [   f       ����                                                                                                                                                                                                                                                                                                                            d   *       d          v       f(�     �   e   f          (                            done <= '0';5��    e                      K
      )               5�_�   [   ]           \   d        ����                                                                                                                                                                                                                                                                                                                            d   *       d          v       f(�     �   c   e   �    �   d   e   �    5��    c                      �	              )       5�_�   \   ^           ]   d       ����                                                                                                                                                                                                                                                                                                                            e   *       e          v       f(�     �   c   e   �      (                            done <= '0';5��    c                     
                     5�_�   ]   _           ^   d       ����                                                                                                                                                                                                                                                                                                                            e   *       e          v       f(�     �   d   f   �    5��    d                      
                     �    d                      
                     5�_�   ^   `           _   Z       ����                                                                                                                                                                                                                                                                                                                            f   *       f          v       f(�     �   Y   [   �                      done <= '1';5��    Y                    	                    5�_�   _   a           `   �   )    ����                                                                                                                                                                                                                                                                                                                            f   *       f          v       f(�8    �   �   �   �      ,                                done <= '1';5��    �   )                 �                    5�_�   `   e           a   ~       ����                                                                                                                                                                                                                                                                                                                            f   *       f          v       f(��     �   }   ~          (                            done <= '1';5��    }                      �      )               5�_�   a   f   b       e   �   )    ����                                                                                                                                                                                                                                                                                                                            f   *       f          v       f(�     �   �   �          ,                                done <= '0';5��    �                      c      -               5�_�   e   g           f   �        ����                                                                                                                                                                                                                                                                                                                            f   *       f          v       f(�	     �   �   �          ,                                done <= '0';5��    �                      G      -               5�_�   f   h           g   �        ����                                                                                                                                                                                                                                                                                                                            f   *       f          v       f(�     �   �   �   �                                  �   �   �   �    5��    �                      �                     �    �                  	                 	       �    �   $                                       5�_�   g   i           h   �   $    ����                                                                                                                                                                                                                                                                                                                            f   *       f          v       f(�     �   �   �   �      $                            done <= 5��    �   $                                       5�_�   h   j           i   �   %    ����                                                                                                                                                                                                                                                                                                                            f   *       f          v       f(�     �   �   �   �      &                            done <= ''5��    �   %                                       5�_�   i   l           j   �   '    ����                                                                                                                                                                                                                                                                                                                            f   *       f          v       f(�     �   �   �   �      '                            done <= '1'5��    �   '                  !                     5�_�   j   m   k       l   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        f(��     �   �   �          5                            if serial_data = '0' then   2                                state <= starting;       *                                -- Control   4                                start_signal <= '1';   2                                shift_data <= '1';                                else5��    �                      #                    5�_�   l   n           m   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        f(��     �   �   �          #                            end if;5��    �                            $               5�_�   m               n   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   f(��   	 �   �   �   �      .                                state <= idle;5��    �                     ?                     5�_�   j           l   k   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f(��     �   �   �        5��    �                      #                    5�_�   a   c       e   b   �   )    ����                                                                                                                                                                                                                                                                                                                            f   *       f          v       f(��     �   �   �   �      ,                                done <= '1';5��    �   )                 �                    5�_�   b   d           c   �   )    ����                                                                                                                                                                                                                                                                                                                            f   *       f          v       f(��     �   �   �   �      ,                                done <= '1';5��    �   )                 �                    5�_�   c               d   �   )    ����                                                                                                                                                                                                                                                                                                                            f   *       f          v       f(��     �   �   �        5��    �                      t      -               5�_�   T   Y   U   [   X   f       ����                                                                                                                                                                                                                                                                                                                            d   *       d          v       f(�     �   e   g        5��    e                      K
      )               5�_�   X   Z           Y   b        ����                                                                                                                                                                                                                                                                                                                            e   *       e          v       f(�     �   b   c   �    �   a   b   �      (                            done <= '0';5��    a                      �	              )       5�_�   Y               Z   b       ����                                                                                                                                                                                                                                                                                                                            e   *       e          v       f(�     �   a   c   �                           done <= '0';5��    a                     �	                     5�_�   T   V       X   U   	       ����                                                                                                                                                                                                                                                                                                                                                             f(�     �      
   �      1        clock, reset, start, serial_data: in bit;5��                         �                      5�_�   U   W           V   d       ����                                                                                                                                                                                                                                                                                                                                                             f(�     �   c   e   �      A                        if start = '1' and serial_data = '0' then5��    c                     
                     5�_�   V               W   �       ����                                                                                                                                                                                                                                                                                                                            d   *       d          v       f(�    �   �   �   �    �   �   �   �      E                            if start = '1' and serial_data = '0' then5��    �                     \                     5�_�   I   K       M   J           ����                                                                                                                                                                                                                                                                                                                            8           9           V        f(�
     �      
        5��                          �       >               5�_�   J   L           K           ����                                                                                                                                                                                                                                                                                                                            7           8           V        f(�     �              5��                          J       #               5�_�   K               L          ����                                                                                                                                                                                                                                                                                                                            7           8           V        f(�     �         �              WIDTH: natural := 75��                         e                      5�_�   F           H   G   I       ����                                                                                                                                                                                                                                                                                                                                                             f(mK     �   H   J   �          clocking: slow_clk5��    H                     	                     �    H                     	                     �    H                                          5�_�   ?           A   @   +       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   *   ,   �      	 )  5��    *                    '                    5�_�   -   /       1   .   �        ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   �   �        5��    �                      �      1               5�_�   .   0           /   �       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   �   �   �       �   �   �   �          end process;5��    �                      �                     �    �                     �                     5�_�   /               0   �       ����                                                                                                                                                                                                                                                                                                                                                  V        f(=�     �   �   �   �          end process;5��    �                     �                     5��