Vim�UnDo� �;B���������qL=����w���8�Gg'   �              e         0       0   0   0    f��    _�       &                      ����                                                                                                                                                                                                                                                                                                                                                             fNE    �   �   �                  wai�   �   �        �       �           �              5��                    �                      �      �    �              '      �              O      5�_�      (          &   I        ����                                                                                                                                                                                                                                                                                                                            I          S          V       f�X    �   H   I                  wait for SERIAL_PERIOD;           serial_data <= '1';            wait for SERIAL_PERIOD;           serial_data <= '1';            wait for SERIAL_PERIOD;           serial_data <= '1';            wait for SERIAL_PERIOD;           serial_data <= '1';            wait for SERIAL_PERIOD;           serial_data <= '1';            wait for SERIAL_PERIOD;5��    H                      ^      Q              5�_�   &   )   '       (   a       ����                                                                                                                                                                                                                                                                                                                            I          I          V       f��     �   a   c   �              �   a   c   �    5��    a                      @	              	       �    a                     H	                     �    a   
                  J	                     �    a   	                  I	                     �    a                    H	                    �    a                    H	                    �    a                 	   H	             	       5�_�   (   *           )   b       ����                                                                                                                                                                                                                                                                                                                            I          I          V       f��     �   a   c   �              reset <= 5��    a                     Q	                     5�_�   )   +           *   b       ����                                                                                                                                                                                                                                                                                                                            I          I          V       f��     �   a   c   �              reset <= ''5��    a                     R	                     5�_�   *   ,           +   b       ����                                                                                                                                                                                                                                                                                                                            I          I          V       f��     �   a   c   �              reset <= '1'5��    a                     T	                     5�_�   +   -           ,   c        ����                                                                                                                                                                                                                                                                                                                            c          o          V       f��     �   b   c                  serial_data <= '1';           wait for SERIAL_PERIOD;           serial_data <= '1';           wait for SERIAL_PERIOD;           serial_data <= '1';      		wait for SERIAL_PERIOD;           serial_data <= '1';           wait for SERIAL_PERIOD;           serial_data <= '1';      		wait for SERIAL_PERIOD;           serial_data <= '1';           wait for SERIAL_PERIOD;           serial_data <= '1';5��    b                      V	      ~              5�_�   ,   .           -   d       ����                                                                                                                                                                                                                                                                                                                            c          c          V       f��     �   d   f   �              �   d   f   �    5��    d                      �	              	       �    d                     �	                     �    d   
                  �	                     �    d   	                  �	                     �    d                    �	                    �    d                    �	                    �    d                 	   �	             	       5�_�   -   /           .   e       ����                                                                                                                                                                                                                                                                                                                            c          c          V       f��     �   d   f   �              reset <= 5��    d                     �	                     5�_�   .   0           /   e       ����                                                                                                                                                                                                                                                                                                                            c          c          V       f��     �   d   f   �              reset <= ''5��    d                     �	                     5�_�   /               0   e       ����                                                                                                                                                                                                                                                                                                                            c          c          V       f��    �   d   f   �              reset <= '0'5��    d                     �	                     5�_�   &           (   '   `       ����                                                                                                                                                                                                                                                                                                                            I          I          V       f��     �   `   a   �       5��    `                      #	              	       �    `                      #	                     5�_�             &      +       ����                                                                                                                                                                                                                                                                                                                                                             fN[    �   *   ,   �      !        while now < 5000 ns loop 5��    *                                        5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             fƫ     �   �   �   �       5��    �                                    	       �    �                                           5�_�                    �        ����                                                                                                                                                                                                                                                                                                                                                             fƯ     �   �   �   �    �   �   �   �              wait for SERIAL_PERIOD;5��    �                                            5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             fƴ     �   �   �   �      "        wait for SERIAL_PERIOD*16;5��    �                     8                     �    �                    9                    5�_�                    �   !    ����                                                                                                                                                                                                                                                                                                                                                             fƻ     �   �   �   �      "        wait for SERIAL_PERIOD*10;5��    �                     :                    5�_�                    �        ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �              �   �   �   �                  reset�   �   �   �              reset <= 5��    �                      =              	       �    �                      =                     �    �                     =              	       �    �                     F                     �    �   	                  G                     �    �                    F                    �    �                    F                    �    �                 
   F             
       �    �                     O                     5�_�      	              �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �              reset <= ''5��    �                     O                     5�_�      
           	   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �              reset <= '1'5��    �                     P                     5�_�   	              
   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �              reset <= '1';5��    �                     R                     5�_�   
                 �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �    �   �   �   �      "        wait for SERIAL_PERIOD*10;5��    �                      T              #       5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      !        wait for SERIAL_PERIOD*4;5��    �                    s                    5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �    �   �   �   �              reset <= '1';5��    �                      v                     5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �              �   �   �   �              start <= 5��    �                      T              	       �    �                     \                     �    �   
                  ^                     �    �   	                  ]                     �    �                    \                    �    �                     `                     �    �                     _                     �    �   
                  ^                     �    �   	                  ]                     �    �                    \                    �    �                    \                    �    �                 	   \             	       5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �              start <= ''5��    �                     e                     5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �              start <= '0'5��    �                     f                     5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �              start <= '0';5��    �                     h                     5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �              reset <= '0';5��    �                    �                    5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �    �   �   �   �      !        wait for SERIAL_PERIOD*4;5��    �                      �              "       5�_�                   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �    �   �   �   �              start <= '0';5��    �                      �                     5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �              start <= '1';5��    �                    �                    5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �              �   �   �   �      	        s5��    �                      �              	       �    �                     �                     5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �    �   �   �   �              start <= '0';5��    �                      �                     5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��    �   �   �        5��    �                      �      
               5�_�                    +       ����                                                                                                                                                                                                                                                                                                                                                             f��    �   *   ,   �      "        while now < 10000 ns loop 5��    *                                        5�_�                    A       ����                                                                                                                                                                                                                                                                                                                                                             f�5     �   @   B   �              wait for 45 ns;5��    @                    �                    5�_�                    A       ����                                                                                                                                                                                                                                                                                                                                                             f�>     �   A   B   �              �   A   C   �              reset <= 5��    A                      �              	       �    A                     �                     �    A   
                  �                     �    A   	                  �                     �    A                    �                    �    A                    �                    �    A                 
   �             
       �    A                     �                     5�_�                    B       ����                                                                                                                                                                                                                                                                                                                                                             f�D     �   A   C   �              reset <= ''5��    A                     �                     5�_�                     B       ����                                                                                                                                                                                                                                                                                                                                                             f�D     �   A   C   �              reset <= '1'5��    A                     �                     5�_�      !               B       ����                                                                                                                                                                                                                                                                                                                                                             f�E     �   A   C   �              reset <= '1';    5��    A                     �                     �    A                    �              	       �    B                      �                     5�_�       #           !   B        ����                                                                                                                                                                                                                                                                                                                            A          B          V       f�J     �   B   C   �    �   B   C   �              wait for 45 ns;           reset <= '1';5��    B                      �              .       5�_�   !   $   "       #   B       ����                                                                                                                                                                                                                                                                                                                            A          B          V       f�U     �   A   C   �              reset <= '0';5��    A                    �                    5�_�   #   %           $   D       ����                                                                                                                                                                                                                                                                                                                            A          B          V       f�V     �   C   E        5��    C                      �                     5�_�   $               %          ����                                                                                                                                                                                                                                                                                                                            A          B          V       f�_    �         �          signal reset : bit := '1';5��                        )                    5�_�   !           #   "   B       ����                                                                                                                                                                                                                                                                                                                            A          B          V       f�O     �   A   C        5��    A                      �                     5�_�                   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �    �   �   �   �              start <= '0';5��    �                      �                     5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �    �   �   �   �      !        wait for SERIAL_PERIOD*4;5��    �                      �              "       5��