Vim�UnDo� '5��R ��C�D�R�}]Q:i�R���N|��   _                                  f(k�    _�                           ����                                                                                                                                                                                                                                                                                                                                                             f(j�     �      	   ^          �      	   ]    5��                          �                      �                          �                      �                        �                     �                     	   �              	       �                         �                      �                         �                      �                        �                     �                         �                      �                         �                      �                     
   �              
       �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �                     
   �              
       �              
          �       
              �                        �                     �                         �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f(j�     �      	   ^          signal not_seg: bit_vector5��                         �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f(j�     �      	   ^           signal not_seg: bit_vector()5��                         �                      �       !                 �                     �       !                 �                     �       !                 �                     5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                                             f(j�     �      	   ^      *    signal not_seg: bit_vector(7 downto 0)5��       *                  �                      5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                             f(j�     �   
      _          �         _    �   
      ^    5��    
                      �                      �    
                     �                     �    
              
       �               �      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f(j�     �         i      .	seg <= 	"1000000" when hex = "0000" else -- 05��                         �                     5�_�      	              %       ����                                                                                                                                                                                                                                                                                                                                                             f(j�     �   &   (   k          seg <= not_seg�   %   (   j          �   %   '   i    5��    %                      8                     �    %                     8                    �    %                      8                     �    %                     8                     �    &                     =                     �    &   	                 B                    �    &                     E                     �    &                    D                    �    &                     F                     �    &                     E                     �    &                    D                    �    &                     J                     �    &                     I                     �    &                     H                     �    &                     G                     �    &                     F                     �    &                     E                     �    &                    D                    �    &                    D                    �    &                    D                    �    &                     J                     �    &                     I                     �    &                     H                     �    &                     G                     �    &                     F                     �    &                     E                     �    &                    D                    �    &                    G                    �    &                     I                     �    &                    H                    �    &                    H                    �    &                    H                    5�_�      
           	   '       ����                                                                                                                                                                                                                                                                                                                                                             f(j�     �   &   (   k          seg <= not not_seg5��    &                     O                     5�_�   	              
   '       ����                                                                                                                                                                                                                                                                                                                                                             f(j�     �   &   (   k          seg <= not not_seg()5��    &                     P                     �    &                    R                    �    &                    R                    �    &                    R                    5�_�   
                 '   "    ����                                                                                                                                                                                                                                                                                                                                                             f(j�     �   &   (   k      $    seg <= not not_seg(6 downto 0)ç   				�   &   (   k      "    seg <= not not_seg(6 downto 0)5��    &   "                  [                     �    &   $                  ]                     �    &   "                 [                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       f(k%     �   
      j      ,            "00111111" when "00110000", -- 05��    
                     �                      �    
   
                  �                      �    
   	                  �                      �    
                     �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       f(k9     �      !   j      )	not_seg <= 	 when hex = "0000" else -- 0    				 when hex = "0001" else -- 1    				 when hex = "0010" else -- 2    				 when hex = "0011" else -- 3    				 when hex = "0100" else -- 4    				 when hex = "0101" else -- 5    				 when hex = "0110" else -- 6    				 when hex = "0111" else -- 7    				 when hex = "1000" else -- 8    				 when hex = "1001" else -- 9   )				"0001000" when hex = "1010" else -- A�         j    �          j   
   2	not_seg <= 	"1000000" when hex = "0000" else -- 0   )				"1001111" when hex = "0001" else -- 1   )				"0100100" when hex = "0010" else -- 2   )				"0110000" when hex = "0011" else -- 3   )				"0011001" when hex = "0100" else -- 4   )				"0010010" when hex = "0101" else -- 5   )				"0000010" when hex = "0110" else -- 6   )				"1111000" when hex = "0111" else -- 7   )				"0000000" when hex = "1000" else -- 8   )				"0010000" when hex = "1001" else -- 95��              	           �      	               �              	           �      	               �              	           �      	               �              	           �      	               �              	                 	               �              	           =      	               �              	           ^      	               �              	                 	               �              	           �      	               �              	           �      	               �                      
   �              
       �                      
   �              
       �                      
   �              
       �                      
                 
       �                      
   D              
       �                      
   o              
       �                      
   �              
       �                      
   �              
       �                      
   �              
       �                      
                 
       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       f(kK     �         k              �         k    �         j    5��                          �              	       �                         �              �       5�_�                           ����                                                                                                                                                                                                                                                                                                                                      &                 f(kQ     �         q      0                "01110111" when "01000001", -- A5��                         �                     5�_�                    '       ����                                                                                                                                                                                                                                                                                                                            '          ,                 f(kx     �   &   .   q       				 when hex = "1010" else -- A    				 when hex = "1011" else -- B    				 when hex = "1100" else -- C    				 when hex = "1101" else -- d    				 when hex = "1110" else -- E    				 when hex = "1111";     -- F    �   '   (   q    �   &   -   q      )				"0001000" when hex = "1010" else -- A   )				"0000011" when hex = "1011" else -- B   )				"1000110" when hex = "1100" else -- C   )				"0100001" when hex = "1101" else -- d   )				"0000110" when hex = "1110" else -- E   )				"0001110" when hex = "1111";     -- F5��    &          	           =      	               �    '          	           ^      	               �    (          	                 	               �    )          	           �      	               �    *          	           �      	               �    +          	           �      	               �    &                  
   =              
       �    '                  
   h              
       �    (                  
   �              
       �    )                  
   �              
       �    *                  
   �              
       �    +                  
                 
       5�_�                   
        ����                                                                                                                                                                                                                                                                                                                            '          ,                 f(k�     �   	   
          			---"gfedcba"5��    	                      �                      5�_�                    
        ����                                                                                                                                                                                                                                                                                                                            &          +                 f(k�     �   	      p    5��    	                      �               	       �    	                     �                     �    	                      �                      5�_�                             ����                                                                                                                                                                                                                                                                                                                            '          ,                 f(k�    �   
             (        "00111111" when "00110000", -- 0   (        "00000110" when "00110001", -- 1   (        "01011011" when "00110010", -- 2   (        "01001111" when "00110011", -- 3   (        "01100110" when "00110100", -- 4   (        "01101101" when "00110101", -- 5   (        "01111101" when "00110110", -- 6   (        "00000111" when "00110111", -- 7   (        "01111111" when "00111000", -- 8   (        "01101111" when "00111001", -- 9   (        "01110111" when "01000001", -- A   (        "01111100" when "01000010", -- B   (        "00111001" when "01000011", -- C   (        "01011110" when "01000100", -- D   (        "01111001" when "01000101", -- E   (        "01110001" when "01000110", -- F        5��    
                      �       �              5�_�                            ����                                                                                                                                                                                                                                                                                                                                                       f(kz     �              5��                          �       �              5�_�                     
        ����                                                                                                                                                                                                                                                                                                                                                             f(i�     �   
      ]                  �         ^    �   
      ^      4                    "00111111" when "00110000", -- 0    5��    
                      �                      �    
                     �                     �    
                     �               )       5��