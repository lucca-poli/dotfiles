Vim�UnDo� �SH\댼�.mKn��1Qd������O&�-=�  W   entity serial_inv is                            f�   
 _�                             ����                                                                                                                                                                                                                                                                                                                                                             f]    �  V              end architecture;�  W            �   �              '            dado_registrado(WIDTH) <= d�   �            �                   �               5��                    �   '                   �      �    �   '           �      �              �      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�     �        W      entity serial_in is5��                         p                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�     �        W      end serial_in;5��              	          �      	              5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�"    �        W      !architecture arch of serial_in is5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�T     �        W      entity serial_in_V0 is5��                         p                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�U     �        W      entity serial_inis5��                         p                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�Z     �        W      $architecture arch of serial_in_V0 is5��                         �                     5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                             f�\    �        W       architecture arch of serial_inis5��                         �                     5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                             f�q     �        W      !architecture arch of serial_in is5��                         �                     5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                             f�w    �        W      entity serial_in is5��                         p                      5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                             f�~     �        W      entity serial_in_ is5��                        p                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f܅    �        W      "architecture arch of serial_in_ is5��                        �                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�O    �        W      entity serial_inV is5��                         p                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f��    �        W      "architecture arch of serial_inV is5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�n     �        W      entity serial_in is5��                         p                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�r   
 �        W      !architecture arch of serial_in is5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�     �        W      !architecture arch of serial_in is5��                         �                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f�	   	 �        W      entity serial_in is5��                         p                      5��