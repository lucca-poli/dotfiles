Vim�UnDo� ��s�"�~�v�2�S	R��`�q����g4�0              	      $       $   $   $    e�L    _�                             ����                                                                                                                                                                                                                                                                                                                                                             e�G�     �                 use IEEE.numeric_std.all;�                   5��                                                  �                                                �                                                �                                                �                                                �                                                �                                                �                                                �                                                �                                                �                                                �                                                �                                                  �                                          D       �                          D                       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�G�     �                 library IEEE;5��                                                  5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�G�     �                 use IEEE.std_logic_1164.all;5��                                                  5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�G�     �                 use IEEE.numeric_std.all;5��                                                5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             e�H
     �                 end entity �                
entity  is�                         �                   5��                                                  �                                                �                                                �                                                �                                                �                                                �                                               �                                                 �                                              �                         1                      �                                                �                         3                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       e�H     �                       5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       e�H     �              5��                                                  5�_�      	                      ����                                                                                                                                                                                                                                                                                                                                                v       e�H     �         	      use IEEE.numeric_std.all;�                 �              5��                                                  �                                                  �                                                �                                                �                                                �                                                �                                                �                                                  �                                          D       �                          D                       5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                v       e�H!     �         	              x, y, z: bit_ve5��                         u                      5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                v       e�H%     �         	              x, y, z: bit_vector5��                         y                      5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                v       e�H&     �         	              x, y, z: bit_vector()5��                         z                      �                        {                     �                        }                     �                        }                     �                        }                     �                        }                     �       1                  �                      �       0                  �                      �       /                  �                      �       .                  �                      �       -                  �                      �       ,                  �                      �       +                  �                      �       *                  �                      �       )                  �                      �       (                  �                      �       '                  �                      �       &                  �                      �       %                  �                      �       $                  �                      �       #                  �                      �       "                  �                      �       !                                        �                          ~                      �                         }                      �                        |                     �       %                  �                      �       $                  �                      �       #                 �                     5�_�                       (    ����                                                                                                                                                                                                                                                                                                                                                v       e�H3     �         	      (        x, y, z: bit_vector(31 downto 0)5��       (                  �                      �       (                 �                     5�_�                       (    ����                                                                                                                                                                                                                                                                                                                                                v       e�H4     �      	   	    �         	    5��                          �               *       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       e�H?     �      	   
      )        x, y, z: bit_vector(31 downto 0);5��                        �                     5�_�                       #    ����                                                                                                                                                                                                                                                                                                                                                v       e�HF     �      	   
      #        q: bit_vector(31 downto 0);5��       "                  �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       e�HI     �      	   
      "        q: bit_vector(31 downto 0)5��                         �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       e�HK    �         
      )        x, y, z: bit_vector(31 downto 0);5��                         o                      5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                v       e�HX     �                 end architecture �               architecture rtl of  is�                     �                 arch�   
               �   
            5��    
                      �                      �    
                      �                      �                          �                      �                         �                      �                         �                      �                         �                      �                         �                     �                         �                     �                         �                     �                         �                     �                        �                      �                          �                       �                        �                      �                                              �                         �                      �                                              5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       e�H_     �             �                 end architecture rtl;�             �             �             �             �             �             �             �             �             �               architecture rtl of ch is5��                        �                     �                                            �                         �                      �                                            �                         �                      �                                            �                         �                      �                                            �                         �                      �                                            �                         �                      �                                            �                         �                      �                                            �                         �                      �                                            �                         �                      �                     	                	       �                         �                      �              	       
         	       
       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       e�H�    �                   5��                         �                      5�_�                      	    ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �                   q <= x or y or z;5��       	                                       5�_�                       	    ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �               
    q <= ;5��       	                                       5�_�                       
    ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �                   q <= ();5��       
                                       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �                   q <= (x and y);5��                                              5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �                   q <= (x and y) xor ;5��                                              5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �                   q <= (x and y) xor ();5��                                              5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �               %    q <= (x and y) xor (not x and y);5��                                              5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �               &    q <= (x and y) xor ((not x and y);5��                         �       '       (       5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �               '    q <= (x and y) xor ((not) x and y);5��                                              5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                                             e�K�     �               &    q <= (x and y) xor ((not x and y);�             5��                                              5�_�       "           !      $    ����                                                                                                                                                                                                                                                                                                                                                             e�L     �               '    q <= (x and y) xor ((not x) and y);5��       $                                     5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                                                             e�L     �                    5��                          �                      5�_�   "   $           #          ����                                                                                                                                                                                                                                                                                                                                                             e�L	    �                    5��                                               5�_�   #               $           ����                                                                                                                                                                                                                                                                                                                                                             e�L    �                 library IEEE;   use IEEE.std_logic_1164.all;   use IEEE.numeric_std.all;    5��                                   F               5�_�                      ,    ����                                                                                                                                                                                                                                                                                                                                                             e�J�     �               +        x, y, z: in bit_vector(31 downto 0)5��       +                  �                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             e�J�     �              5��                          S                      5��