Vim�UnDo� N��P��;Dh𨟪t$�~}[O_�V�D2�   �   !            assert serial_o = '1'   �                           fA�    _�                            ����                                                                                                                                                                                                                                                                                                                                                             f�Y     �         �      end serial_out_tb;5��                                               5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f�[    �          �      entity serial_out_tb is   end;�         �      end;5��                                                �                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                      &           V       fȁ    �                    component serial_out2       generic (   $        POLARITY  : boolean := TRUE;   !        WIDTH     : natural := 8;   !        PARITY    : natural := 1;            STOP_BITS : natural := 1       );   
    port (           clock    : in  bit;           reset    : in  bit;           tx_go    : in  bit;           tx_done  : out bit;   4        data     : in  bit_vector(WIDTH-1 downto 0);           serial_o : out bit       );       end component;    5��                          "      �              5�_�                     �        ����                                                                                                                                                                                                                                                                                                                                                             fA�    �   �   �   �      !            assert serial_o = '1'5��    �                      �                     �    �                      �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�f     �         �          component serial_out5��                         :                     5��