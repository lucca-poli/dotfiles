Vim�UnDo� Z��8TOuW�L�m�5�Ȣ8)���s��Ǻ�   ]   \    out_multisteps: multisteps port map (CLOCK_50, not KEY(1), generic_in, result, LEDR(0));   R   )                       f��    _�                             ����                                                                                                                                                                                                                                                                                                                                       o           V        f�    �                  entity interface is�               �             n   
    port (   +        input : in bit_vector (7 downto 0);   .        selected : in bit_vector (1 downto 0);   -        result : out bit_vector (31 downto 0)       );   end interface;       *architecture arc_interface of interface is       component stepfun is   		port (   >			ai, bi, ci, di, ei, fi, gi, hi: in bit_vector(31 downto 0);   #			kpw: in bit_vector(31 downto 0);   >			ao, bo, co, do, eo, fo, go, ho: out bit_vector(31 downto 0)   		);       end component;       1    signal generic_in : bit_vector (31 downto 0);   E    signal ao, bo, co, do, eo, fo, go, ho : bit_vector (31 downto 0);       begin   0    generic_in <= input & input & input & input;       �    out_stepfun: stepfun port map (generic_in, generic_in, generic_in, generic_in, generic_in, generic_in, generic_in, generic_in, generic_in, ao, bo, co, do, eo, fo, go, ho);       ,    result <= ao when (selected = "01") else    		eo when (selected = "10") else   		bo;       end arc_interface;       entity hex2seg is   ,    port ( hex : in  bit_vector(3 downto 0);   +           seg : out bit_vector(6 downto 0)   
        );   end hex2seg;       )architecture comportamental of hex2seg is   begin   			---"gfedcba"   .	seg <= 	"1000000" when hex = "0000" else -- 0   )				"1001111" when hex = "0001" else -- 1   )				"0100100" when hex = "0010" else -- 2   )				"0110000" when hex = "0011" else -- 3   )				"0011001" when hex = "0100" else -- 4   )				"0010010" when hex = "0101" else -- 5   )				"0000010" when hex = "0110" else -- 6   )				"1111000" when hex = "0111" else -- 7   )				"0000000" when hex = "1000" else -- 8   )				"0010000" when hex = "1001" else -- 9   )				"0001000" when hex = "1010" else -- A   )				"0000011" when hex = "1011" else -- B   )				"1000110" when hex = "1100" else -- C   )				"0100001" when hex = "1101" else -- d   )				"0000110" when hex = "1110" else -- E   )				"0001110" when hex = "1111";     -- F   				       end comportamental;           entity board is   	    port(   '        SW : in bit_vector(9 downto 0);       )        HEX0: out bit_vector(6 downto 0);   )        HEX1: out bit_vector(6 downto 0);   )        HEX2: out bit_vector(6 downto 0);   )        HEX3: out bit_vector(6 downto 0);   )        HEX4: out bit_vector(6 downto 0);   )        HEX5: out bit_vector(6 downto 0);       (        LEDR: out bit_vector(9 downto 0)       );   
end board;       #architecture behavioral of board is   4    signal selected_output : bit_vector(1 downto 0);   (	 signal sinal : bit_vector(7 downto 0);   +    signal result: bit_vector(31 downto 0);               component hex2seg is    -        port (hex: in bit_vector(3 downto 0);   +            seg: out bit_vector(6 downto 0)               );       end component;           component interface is   
    port (   +        input : in bit_vector (7 downto 0);   .        selected : in bit_vector (1 downto 0);   -        result : out bit_vector (31 downto 0)       );       end component;   begin   &    selected_output <= SW(9 downto 8);   	 sinal <= SW(7 downto 0);   d	 interface_comp: interface port map(input => sinal, selected => selected_output, result => result);       I    HEX0_comp: hex2seg port map (hex => result(3 downto 0), seg => HEX0);   I    HEX1_comp: hex2seg port map (hex => result(7 downto 4), seg => HEX1);   J    HEX2_comp: hex2seg port map (hex => result(11 downto 8), seg => HEX2);   K    HEX3_comp: hex2seg port map (hex => result(15 downto 12), seg => HEX3);   K    HEX4_comp: hex2seg port map (hex => result(19 downto 16), seg => HEX4);   K    HEX5_comp: hex2seg port map (hex => result(23 downto 20), seg => HEX5);   	    2	 LEDR(9 downto 8) <= "00"; -- Leds 8 e 9 apagados   -    LEDR(7 downto 0) <= result(31 downto 24);   	    end architecture;5��           n                      y              �                                                  �                    i                      �      5�_�                            ����                                                                                                                                                                                                                                                                                                                                       j           V        f��     �                  entity interface is�               �             i   
    port (   +        input : in bit_vector (7 downto 0);   		  rst, clk: in bit;   		  done: out bit;   .        result : out bit_vector (255 downto 0)       );   end interface;       *architecture arc_interface of interface is       component multisteps is   		port (   		  clk, rst : in bit;   +        msgi : in bit_vector(511 downto 0);   ,        haso : out bit_vector(255 downto 0);           done : out bit   		);       end component;       2    signal generic_in : bit_vector (511 downto 0);       begin      generic_in <= input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input;       M    out_multisteps: multisteps port map (clk, rst, generic_in, result, done);       end arc_interface;       entity hex2seg is   ,    port ( hex : in  bit_vector(3 downto 0);   +           seg : out bit_vector(6 downto 0)   
        );   end hex2seg;       )architecture comportamental of hex2seg is   begin   			---"gfedcba"   .	seg <= 	"1000000" when hex = "0000" else -- 0   )				"1001111" when hex = "0001" else -- 1   )				"0100100" when hex = "0010" else -- 2   )				"0110000" when hex = "0011" else -- 3   )				"0011001" when hex = "0100" else -- 4   )				"0010010" when hex = "0101" else -- 5   )				"0000010" when hex = "0110" else -- 6   )				"1111000" when hex = "0111" else -- 7   )				"0000000" when hex = "1000" else -- 8   )				"0010000" when hex = "1001" else -- 9   )				"0001000" when hex = "1010" else -- A   )				"0000011" when hex = "1011" else -- B   )				"1000110" when hex = "1100" else -- C   )				"0100001" when hex = "1101" else -- d   )				"0000110" when hex = "1110" else -- E   )				"0001110" when hex = "1111";     -- F   				       end comportamental;           entity board is   	    port(   '        SW : in bit_vector(9 downto 0);   #		  KEY: in bit_vector(9 downto 0);   		  CLK: in bit;       )        HEX0: out bit_vector(6 downto 0);   )        HEX1: out bit_vector(6 downto 0);   )        HEX2: out bit_vector(6 downto 0);   )        HEX3: out bit_vector(6 downto 0);   )        HEX4: out bit_vector(6 downto 0);   )        HEX5: out bit_vector(6 downto 0);       (        LEDR: out bit_vector(9 downto 0)       );   
end board;       #architecture behavioral of board is   ,    signal result: bit_vector(255 downto 0);           component hex2seg is    -        port (hex: in bit_vector(3 downto 0);   +            seg: out bit_vector(6 downto 0)               );       end component;           component interface is   
    port (   +        input : in bit_vector (7 downto 0);   		  rst, clk: in bit;   		  done: out bit;   .        result : out bit_vector (255 downto 0)       );       end component;   begin       W	 interface_comp: interface port map(SW(7 downto 0), not KEY(1), CLK, LEDR(0), result);       I    HEX0_comp: hex2seg port map (hex => result(3 downto 0), seg => HEX0);   I    HEX1_comp: hex2seg port map (hex => result(7 downto 4), seg => HEX1);   J    HEX2_comp: hex2seg port map (hex => result(11 downto 8), seg => HEX2);   K    HEX3_comp: hex2seg port map (hex => result(15 downto 12), seg => HEX3);   K    HEX4_comp: hex2seg port map (hex => result(19 downto 16), seg => HEX4);   K    HEX5_comp: hex2seg port map (hex => result(23 downto 20), seg => HEX5);   	    	 LEDR(1) <= not KEY(1);   	    end architecture;5��           i                      |              �                                                  �                    R                      �      5�_�                   2        ����                                                                                                                                                                                                                                                                                                                            2          6          V       f��     �   1   7   S          component hex2seg is    -        port (hex: in bit_vector(3 downto 0);   +            seg: out bit_vector(6 downto 0)               );       end component;5�5�_�                   1        ����                                                                                                                                                                                                                                                                                                                            2           6           V        f�     �   0   2   S    5��    0                      _                     �    0                      _                     �    0                      _                     5�_�      	              1        ����                                                                                                                                                                                                                                                                                                                            3           7           V        f�     �   1   7   T    �   1   2   T    5��    1                      `              �       5�_�      
           	   2       ����                                                                                                                                                                                                                                                                                                                            8           <           V        f�
     �   1   3   Y          component hex2seg is 5��    1                    n                    �    1                     p                     �    1                     o                     �    1                    n                    5�_�   	              
   3       ����                                                                                                                                                                                                                                                                                                                            3          4   +       v���    f�     �   3   6   X    �   2   5   W              port (            );�   3   4   W    �   2   4   Y      -        port (hex: in bit_vector(3 downto 0);   +            seg: out bit_vector(6 downto 0)               );5��    2                     �      L               �    2                     �              2       5�_�   
                 4       ����                                                                                                                                                                                                                                                                                                                            4           5          v���    f�      �   3   5   Z              clk_in: in bit;5��    3                     �                     5�_�                    5       ����                                                                                                                                                                                                                                                                                                                            4           5          v���    f�!    �   4   6   Z              clk_out: out bit5��    4                     �                     5�_�                    O        ����                                                                                                                                                                                                                                                                                                                                                             f�]     �   N   P   [          �   N   P   Z    5��    N                      �	                     �    N                     �	                     �    N                     
                     �    N                      
                     �    N                     �	                     �    N                     �	                     �    N   
                  �	                     �    N   	                  �	                     �    N                     �	                     �    N                    �	                    �    N                     
                     �    N                      
                     �    N                    �	                    �    N                    �	                    �    N                    �	                    �    N                     

                     �    N                     	
                     �    N                    
                    �    N                    
                    �    N                 	   
             	       5�_�                    O       ����                                                                                                                                                                                                                                                                                                                                                             f�o     �   N   P   [          clking: slow_clk port map 5��    N                     
                     5�_�                    O       ����                                                                                                                                                                                                                                                                                                                                                             f�p     �   N   P   [           clking: slow_clk port map ()5��    N                     
                     �    N                    
                    �    N                    
                    �    N                 
   
             
       5�_�                    B       ����                                                                                                                                                                                                                                                                                                                            B          D                 f�}     �   B   E   [      ,        haso : out bit_vector(255 downto 0);           done : out bit�   A   C   [      +        msgi : in bit_vector(511 downto 0);5��    A                     �                     �    B                     �                     �    C                     "                     5�_�                    A       ����                                                                                                                                                                                                                                                                                                                            B          D                 f�     �   @   B   [      		  clk, rst : in bit;5��    @                     �                     5�_�                    :       ����                                                                                                                                                                                                                                                                                                                            B          D                 f��     �   9   <   [      -        port (hex: in bit_vector(3 downto 0);5��    9                                  	       �    :                                         5�_�                    ;       ����                                                                                                                                                                                                                                                                                                                            C          E                 f��     �   :   <   \      0                 hex: in bit_vector(3 downto 0);5��    :                                          5�_�                    ;       ����                                                                                                                                                                                                                                                                                                                            C          E                 f��     �   :   <   \      /                hex: in bit_vector(3 downto 0);5��    :                                          5�_�                    =       ����                                                                                                                                                                                                                                                                                                                            C          E                 f��     �   <   >   \                  );5��    <                     o                     5�_�                    6       ����                                                                                                                                                                                                                                                                                                                            C          E                 f��     �   5   7   \                  );5��    5                     �                     5�_�                   K   	    ����                                                                                                                                                                                                                                                                                                                            C          E                 f��     �   K   M   ]           �   K   M   \    5��    K                      �                     �    K                     �                     �    K                     �                     �    K                     �                     �    K                     �                     �    K                    �                    5�_�                    Q   )    ����                                                                                                                                                                                                                                                                                                                            C          E                 f��     �   P   R   ]      *    clking: slow_clk port map (CLOCK_50, )5��    P   )                  I
                     �    P   )                 I
                    �    P   )                 I
                    �    P   )                 I
                    �    P   )                 I
                    �    P   )                 I
                    5�_�                    Q   1    ����                                                                                                                                                                                                                                                                                                                            C          E                 f��     �   P   R   ]      1    clking: slow_clk port map (CLOCK_50, art_clk)5��    P   1                  Q
                     5�_�                     R   )    ����                                                                                                                                                                                                                                                                                                                            C          E                 f��    �   Q   S   ]      \    out_multisteps: multisteps port map (CLOCK_50, not KEY(1), generic_in, result, LEDR(0));5��    Q   )                 |
                    �    Q   +                  ~
                     �    Q   *                  }
                     �    Q   )                 |
                    �    Q   )                 |
                    �    Q   )                 |
                    5�_�                    K   	    ����                                                                                                                                                                                                                                                                                                                            C          E                 f��     �   J   K   \           �   J   L   ]           u5��    J                      �                     �    J                     �                     5�_�                   1        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   1   2   S    �   1   2   S   j   entity interface is   
    port (   +        input : in bit_vector (7 downto 0);   		  rst, clk: in bit;   		  done: out bit;   .        result : out bit_vector (255 downto 0)       );   end interface;       *architecture arc_interface of interface is       component multisteps is   		port (   		  clk, rst : in bit;   +        msgi : in bit_vector(511 downto 0);   ,        haso : out bit_vector(255 downto 0);           done : out bit   		);       end component;       2    signal generic_in : bit_vector (511 downto 0);       begin      generic_in <= input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input & input;       M    out_multisteps: multisteps port map (clk, rst, generic_in, result, done);       end arc_interface;       entity hex2seg is   ,    port ( hex : in  bit_vector(3 downto 0);   +           seg : out bit_vector(6 downto 0)   
        );   end hex2seg;       )architecture comportamental of hex2seg is   begin   			---"gfedcba"   .	seg <= 	"1000000" when hex = "0000" else -- 0   )				"1001111" when hex = "0001" else -- 1   )				"0100100" when hex = "0010" else -- 2   )				"0110000" when hex = "0011" else -- 3   )				"0011001" when hex = "0100" else -- 4   )				"0010010" when hex = "0101" else -- 5   )				"0000010" when hex = "0110" else -- 6   )				"1111000" when hex = "0111" else -- 7   )				"0000000" when hex = "1000" else -- 8   )				"0010000" when hex = "1001" else -- 9   )				"0001000" when hex = "1010" else -- A   )				"0000011" when hex = "1011" else -- B   )				"1000110" when hex = "1100" else -- C   )				"0100001" when hex = "1101" else -- d   )				"0000110" when hex = "1110" else -- E   )				"0001110" when hex = "1111";     -- F   				       end comportamental;           entity board is   	    port(   '        SW : in bit_vector(9 downto 0);   #		  KEY: in bit_vector(9 downto 0);   		  CLK: in bit;       )        HEX0: out bit_vector(6 downto 0);   )        HEX1: out bit_vector(6 downto 0);   )        HEX2: out bit_vector(6 downto 0);   )        HEX3: out bit_vector(6 downto 0);   )        HEX4: out bit_vector(6 downto 0);   )        HEX5: out bit_vector(6 downto 0);       (        LEDR: out bit_vector(9 downto 0)       );   
end board;       #architecture behavioral of board is   ,    signal result: bit_vector(255 downto 0);           component hex2seg is    -        port (hex: in bit_vector(3 downto 0);   +            seg: out bit_vector(6 downto 0)               );       end component;           component interface is   
    port (   +        input : in bit_vector (7 downto 0);   		  rst, clk: in bit;   		  done: out bit;   .        result : out bit_vector (255 downto 0)       );       end component;   begin       W	 interface_comp: interface port map(SW(7 downto 0), not KEY(1), CLK, LEDR(0), result);       I    HEX0_comp: hex2seg port map (hex => result(3 downto 0), seg => HEX0);   I    HEX1_comp: hex2seg port map (hex => result(7 downto 4), seg => HEX1);   J    HEX2_comp: hex2seg port map (hex => result(11 downto 8), seg => HEX2);   K    HEX3_comp: hex2seg port map (hex => result(15 downto 12), seg => HEX3);   K    HEX4_comp: hex2seg port map (hex => result(19 downto 16), seg => HEX4);   K    HEX5_comp: hex2seg port map (hex => result(23 downto 20), seg => HEX5);   	    	 LEDR(1) <= not KEY(1);   	    end architecture;5��    1               j       `              �      5�_�                    1        ����                                                                                                                                                                                                                                                                                                                            4          8          V       f��     �   0   1   S          �   0   2   T           5��    0                      _                     �    0                      _                     �    0                      _                     �    0                     _                     �    1                      `                     5�_�                    0       ����                                                                                                                                                                                                                                                                                                                                       V           V        f��     �   0   1   S          �   0   2   T           5��    0                      _                     �    0                      _                     �    0                      _                     �    0                     _                     �    1                      `                     5��