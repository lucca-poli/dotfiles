Vim�UnDo� ��s���I�q���2Z��KB�j/'��{�Hh�   S   W        "Did not proceed to 4, count is " & integer'image(to_integer(unsigned(count)))    A   :      0       0   0   0    f�    _�                     	        ����                                                                                                                                                                                                                                                                                                                            	                      V        f��     �         M    �   	   
   M    �      	          C            clk : in bit;                            -- Clock input   A            rst : in bit;                          -- Reset input   F            count : out integer       -- 6-bit count output (64 steps)5��                          �       �               �                          �               �       5�_�                    	       ����                                                                                                                                                                                                                                                                                                                            	                           f��     �   	      P              done: out bit;   B        count : out natural       -- 6-bit count output (64 steps)�      
   P      J        clk, rst, start: in bit;                            -- Clock input5��                         �                      �    	                     �                      �    
                     	                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         P      -    signal rst : bit := '0';  -- Reset signal5��                        �                    �                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         P      -    signal clk : bit := '0';  -- Clock signal5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         P      /    signal clk,  : bit := '0';  -- Clock signal�         P    5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         P      2    signal clk, rst : bit := '0';  -- Clock signal5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f�     �         P      8    signal clk, rst, done : bit := '0';  -- Clock signal5��                         �                     5�_�      	                     ����                                                                                                                                                                                                                                                                                                                            	                           f�     �                *    signal  : bit := '0';  -- Reset signal5��                          �      +               5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                            	                           f�     �         O          component counter_6bit5��                        �                     5�_�   	              
   !   	    ����                                                                                                                                                                                                                                                                                                                            !   	       !          v       f�!     �       "   O          dut: counter_6bit�   !   "   O    5��        	                 H                    5�_�   
                 $        ����                                                                                                                                                                                                                                                                                                                            !   	       !          v       f�*     �   "   $   M                  clk => clk,�   #   $                      rst => rst,               count => count5��    #                      �      3               �    "                     w                     �    "                     k                    �    "                     l                     �    "                      k                     5�_�                    $       ����                                                                                                                                                                                                                                                                                                                            !   	       !          v       f�,     �   !   #   K              port map (clk, rst);�   !   #   L              port map (   );�   "   $   M          );�   #   %   M      
        );5��    #                     m                     �    #                      l                     �    "                      k                     �    !                     j                     �    !                     j                     �    !                     p                     �    !                    o                    �    !                    o                    �    !                    o                    �    !                    t                    �    !                     u                     �    !                    t                    �    !                    t                    �    !                 	   t             	       �    !   $                  |                     �    !   #                 {                    �    !   #                 {                    �    !   #              	   {             	       �    !   +                  �                     �    !   *                  �                     �    !   )                 �                    �    !   )                 �                    �    !   )                 �                    5�_�                    E       ����                                                                                                                                                                                                                                                                                                                            !   	       !          v       f�X     �   E   H   L              �   E   G   K    5��    E                                    	       �    E                                           �    E                                   	       �    F                                           5�_�                    G        ����                                                                                                                                                                                                                                                                                                                            !   	       !          v       f�Y     �   G   I   M    �   G   H   M    5��    G                                           5�_�                    G        ����                                                                                                                                                                                                                                                                                                                            !   	       !          v       f�Z     �   F   G           5��    F                                           5�_�                           ����                                                                                                                                                                                                                                                                                                                            !   	       !          v       f�p     �         M    �         M    5��                          �              @       5�_�                           ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       f�s     �         N      ?    signal clk, rst, start, done : bit := '0';  -- Clock signal5��              
                 
               5�_�                           ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       f�v     �         N      5    signal start, done : bit := '0';  -- Clock signal5��                                              5�_�                           ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       f�y     �         N      .    signal start: bit := '0';  -- Clock signal5��                                            5�_�                           ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       f�|     �         N      ?    signal clk, rst, start, done : bit := '0';  -- Clock signal5��                         �                     5�_�                    1       ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       fҌ     �   0   2   O              �   0   2   N    5��    0                      �              	       �    0                     �                     �    0   
                  �                     �    0   	                  �                     �    0                    �                    �    0                    �                    �    0                 	   �             	       5�_�                    1       ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       fґ     �   0   2   O              start <= 5��    0                     �                     5�_�                    1       ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       fґ     �   0   2   O              start <= ''5��    0                                           5�_�                    1       ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       fғ     �   0   2   O              start <= '0'5��    0                                          5�_�                    #       ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       fҡ     �   "   $   O    �   #   $   O    5��    "                      �              1       5�_�                    #       ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       fҢ     �   "   $   P      0        port map (clk, rst, start, done, count);5��    "                    �                    5�_�                    #       ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       fҩ     �   "   $   P      3        generic map (clk, rst, start, done, count);5��    "                    �                    �    "                    �                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       f��     �         P    �         P    5��                          �               /       5�_�                           ����                                                                                                                                                                                                                                                                                                                                      
                 f��     �         S              MAX_COUNT: natural       );�      	   S          generic(5��                         �                      �                         �                      �    	                     �                      5�_�                    &       ����                                                                                                                                                                                                                                                                                                                                      
                 f��     �   %   '   S              generic map (8);5��    %                     �                     5�_�                     1   E    ����                                                                                                                                                                                                                                                                                                                                      
                 f��     �   0   2   S      V        "Did not proceed to 1, count is " & integer'image(to_integer(unsigned(count)))5��    0   E                  �                     5�_�      !               1   E    ����                                                                                                                                                                                                                                                                                                                                      
                 f��     �   0   2   S      N        "Did not proceed to 1, count is " & integer'image(to_integer((count)))5��    0   E                  �                     5�_�       "           !   1   J    ����                                                                                                                                                                                                                                                                                                                                      
                 f��     �   0   2   S      M        "Did not proceed to 1, count is " & integer'image(to_integer(count)))5��    0   J                  �                     5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                                      
                 f��     �         S      .    signal count : integer;  -- Input stimulus5��                        l                    �                         q                     �                         p                     �                         o                     �                         n                     �                         m                     �                        l                    �                        l                    �                        l                    5�_�   "   $           #   1   :    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   0   2   S      L        "Did not proceed to 1, count is " & integer'image(to_integer(count))5��    0   :       
           �      
               5�_�   #   %           $   1   :    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   0   2   S      B        "Did not proceed to 1, count is " & integer'image((count))5��    0   :                  �                     5�_�   $   &           %   1   ?    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   0   2   S      A        "Did not proceed to 1, count is " & integer'image(count))5��    0   ?                  �                     5�_�   %   '           &   7   :    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   6   8   S      V        "Did not proceed to 2, count is " & integer'image(to_integer(unsigned(count)))5��    6   :                  �                     5�_�   &   (           '   7   9    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   6   8   S      C        "Did not proceed to 2, count is " & integer'image((count)))5��    6   9                  �                     5�_�   '   )           (   7   ?    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   6   8   S      B        "Did not proceed to 2, count is " & integer'image(count)))5��    6   ?                  �                     5�_�   (   *           )   7   ?    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   6   8   S      A        "Did not proceed to 2, count is " & integer'image(count))5��    6   ?                  �                     5�_�   )   +           *   <   :    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   ;   =   S      V        "Did not proceed to 3, count is " & integer'image(to_integer(unsigned(count)))5��    ;   :                  6                     5�_�   *   ,           +   <   :    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   ;   =   S      C        "Did not proceed to 3, count is " & integer'image((count)))5��    ;   :                  6                     5�_�   +   -           ,   <   ?    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   ;   =   S      B        "Did not proceed to 3, count is " & integer'image(count)))5��    ;   ?                  ;                     5�_�   ,   .           -   <   ?    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   ;   =   S      A        "Did not proceed to 3, count is " & integer'image(count))5��    ;   ?                  ;                     5�_�   -   /           .   A   :    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   @   B   S      W        "Did not proceed to 4, count is " & integer'image(to_integer(unsigned(count))) 5��    @   :                  �                     5�_�   .   0           /   A   ?    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   @   B   S      C        "Did not proceed to 4, count is " & integer'image(count))) 5��    @   ?                  �                     5�_�   /               0   A   ?    ����                                                                                                                                                                                                                                                                                                                                      
                 f�    �   @   B   S      B        "Did not proceed to 4, count is " & integer'image(count)) 5��    @   ?                  �                     5��