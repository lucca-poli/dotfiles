Vim�UnDo� �wLK}x��r�SI��c��|�E���| ���(�      -            if counter = (others => '1') then                                 f��    _�                             ����                                                                                                                                                                                                                                                                                                                                                             f��     �                 end entity �                
entity  is�                         �                   5��                                                  �                                                �                                                �                                                �                                                �                                                �                                                �                                               �                                                 �                                              �                         1                      �                                                �                         9                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f��     �                       5��                         &                      �                        4                     �                        5               	       �                         6                     �                        A                     �                        K                     �                         N                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f�     �                 end architecture �      	         architecture rtl of  is�                     �                 arch�                 end entity slow_clk;5��                         j                      �                          k                      �                          l                      �                         n                      �                         m                      �                         l                     �                         l                     �                         l                     �                         l                     �                        �                      �                          �                       �                        �                      �                         �                      �                         �                      �                         �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f�     �      	       �                 end architecture rtl;�      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	       �      	         architecture rtl of slow_clk is5��                        y                     �                        �                     �                         z                      �                        �                     �                         {                      �                        �                     �                         |                      �                        �                     �                         }                      �                        �                     �                         ~                      �                        �                     �                                               �                        �                     �                         �                      �                        �                     �                         �                      �                     	   �              	       �                         �                      �              	       
   �       	       
       �                         �                      �              
       	   �       
       	       �                         �                      �              	          �       	              �                         �                      �                        �                     �                                               �                        �                     �                         ~                      �                        �                     �                         }                      �                        �                     �                         |                      �                        �                     �                         {                      �                        �                     �                         z                      �                        �                     �                         y                      �                         �                      �                         y                      �                         �                      �                         z                      �                        �                     �                         {                      �                        �                     5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                v       f�&     �   	                signal counter: uns�                   �      
       5��                          �                      �                          �                      �                         �                      �    	                     �                      �    	                     �                      �    	                     �                      �    	                    �                     �    	                    �                     �    	                    �                     �    	                    �                     5�_�                    
       ����                                                                                                                                                                                                                                                                                                                            
          
          v       f�G     �   	            (    signal counter: unsigned(7 downto 0)5��    	                    �                     5�_�                    
   (    ����                                                                                                                                                                                                                                                                                                                            
   &       
   &       v   &    f�K     �   	            (    signal counter: unsigned(9 downto 0)5��    	   (                  �                      5�_�      	                     ����                                                                                                                                                                                                                                                                                                                            
   &       
   &       v   &    f�P     �              5��                                                  5�_�      
           	           ����                                                                                                                                                                                                                                                                                                                               &          &       v   &    f�Q     �               use IEEE.numeric_std.all;�                 �              5��                                                  �                                                  �                                                �                                                �                                                �                                                �                                                �                                                  �                                          D       �                          D                       5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                               &          &       v   &    f�T     �                use IEEE.std_logic_1164.all;5��                                                5�_�   
                    	    ����                                                                                                                                                                                                                                                                                                                               &          &       v   &    f�U     �               use IEEE.numeric_std.all;5��       	                                      �                                               �       
                                        �       	                                      �                                               �       
                                        �       	                                      �       	                                      �       	                                      �       	                                      5�_�                           ����                                                                                                                                                                                                                                                                                                                               &          &       v   &    f�[     �                   end process �                       if rising_edge() then�                               �                           if �                       if �                   5��                         �                      �                        �                     �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                                              �                                              �                                               �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                        �                     �                        �                     �                        �                     �                        
                     �                         !                     �                        -                     �                         C                     �                        P                     �                          f                      �                        f              W       �                         �                     �                         -                     �                      	   �              	       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f��     �             �                   end process proc_name;�             �             �             �             �             �                   proc_name: process(clk)5��              	          �       	              �              	          �      	              �                         �                      �                        �                    �                         �                      �                        �                    �                         �                      �                        �                    �                         �                      �                        �                    �       	                  �                      �                        �                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f�     �                   timing: process(clk_in)�             �                        if rising_edge(clk) then�             �             �             �             �             �             �             �             �             �             �             �                   timing: process(clk)5��                                            �                        (                    �                                              �                        )                    �                                              �                        *                    �                                              �                        )                    �                                              �                        (                    �                                              �                         '                     �                                              �                         (                     �                                              �                        )                    �                                              �                        *                    �                                              �                        +                    �                                              �                        ,                    �                         	                     �                        -                    �                         	                     �                                              �                                              �                                              �                                              �                                            �                                            �                                            5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       f�     �                !            if rst = rst_val then                                  else                                  end if;5��                          :      i               5�_�                          ����                                                                                                                                                                                                                                                                                                                                                V       f��     �                       end if;5��                           :                      5�_�                          ����                                                                                                                                                                                                                                                                                                                                                V       f��    �                       end if;5��                           :                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f��     �                               �                           �             5��                          :              	       �                         :                    �                         G                     �                        F                    �                         G                     �                        F                    �                        F                    �                        F                    �                        F                    �                        R                     �                          h                      �                        h                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f��     �                           if condition then5��              	          I      	              �                         L                     �                         K                     �                         J                     �                        I                    �                        I                    �                     
   I             
       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f��     �                           if counter =  then5��                         S                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f��     �                            if counter = () then5��                         T                     �                         V                     �                         U                     �                        T                    �                        T                    �                        T                    �                        T                    5�_�                       &    ����                                                                                                                                                                                                                                                                                                                                                v       f��     �               -            if counter = (others => '0') then5��       %                 _                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f��     �                               5��                         x                     �                         z                     �                         y                     �                        x                    �                         }                     �                         |                     �                         {                     �                         z                     �                         y                     �                        x                    �                         ~                     �                         }                     �                         |                     �                         {                     �                         z                     �                         y                     �                        x                    �                        x                    �                        x                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f��     �                   �             5��                          �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                        �                     �                        �                     �                     	   �              	       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f��     �                               clk_out5��                      
   �              
       �                          �                     �                        �                    �                        �                    �                        �                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f�     �                   signal current_state: bit;5��                         �                      �       "                                       �       !                                     �       !                                     �       !                                     �       !                                     �       !                                     5�_�                       &    ����                                                                                                                                                                                                                                                                                                                                                v       f�%    �                           �             5��                          c                     �                         o                     �                         r                     �                         q                     �                         p                     �                        o                    �                        o                    �                        o                    �                         }                     �                         |                     �                         {                     �                        z                    �                        z                    �                        z                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �               -            if counter = (others => '1') then5��                         �                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �                           if counter =  then5��                         �                     5�_�                             ����                                                                                                                                                                                                                                                                                                                                                  V        f��    �                            if counter = "" then5��                      
   �              
       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       f��     �                �                                                  end if;�             �                                       end if;5��                          :              	       �                         :                    �                         G                     �                         E                     �       
                  D                     �       	                  C                     �                         B                     �                         A                     �                         @                     �                         ?                     �                         >                     �                         =                     �                         <                     �                         ;                     �                          :                     �                       ;                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f�     �                           �               1            generate_label: if condition generate                   �                                              end generate �               (            end generate generate_label;5��                          :              	       �                         :                    �                         H                     �                         G                     �                        F                    �                        F                    �                        F                    �                        F                    �       (                 b                     �                          |                      �                        |                     �                         �                     5��