Vim�UnDo� 5 �&���Q��КC"��$jW��<��η   �                                  f;xi    _�                     o   ,    ����                                                                                                                                                                                                                                                                                                                                                             f;w5     �   n   p   �      /                                tx_done <= '0';5��    n   ,                 �                    5�_�                    X   +    ����                                                                                                                                                                                                                                                                                                                                                             f;w;     �   X   Z   �                              �   X   Z   �    5��    X                      �	                     �    X                     	
                     �    X                     

                     �    X                    	
                    �    X                     
                     �    X                     
                     �    X                     
                     �    X                     

                     �    X                    	
                    �    X                     
                     �    X                     
                     �    X                     
                     �    X                     
                     �    X                     
                     �    X                     

                     �    X                    	
                    �    X                    	
                    �    X                    	
                    5�_�                    Y   #    ����                                                                                                                                                                                                                                                                                                                                                             f;w@     �   X   Z   �      #                        tx_done <= 5��    X   #                  
                     5�_�                    Y   $    ����                                                                                                                                                                                                                                                                                                                                                             f;w@     �   X   Z   �      %                        tx_done <= ''5��    X   $                  
                     5�_�                    Y   &    ����                                                                                                                                                                                                                                                                                                                                                             f;wA    �   X   Z   �      &                        tx_done <= '0'5��    X   &                  
                     5�_�                    b   "    ����                                                                                                                                                                                                                                                                                                                                                             f;x3     �   b   d   �                                  �   b   d   �    5��    b                      �                     �    b                     �                     �    b                     �                     �    b                     �                     �    b                    �                    �    b                    �                    �    b                    �                    5�_�                    c   '    ����                                                                                                                                                                                                                                                                                                                                                             f;x8     �   b   d   �      '                            tx_done <= 5��    b   '                  �                     5�_�      	              c   (    ����                                                                                                                                                                                                                                                                                                                                                             f;x8     �   b   d   �      )                            tx_done <= ''5��    b   '                  �                     �    b   '                  �                     5�_�      
           	   c   '    ����                                                                                                                                                                                                                                                                                                                                                             f;x9     �   b   d   �      '                            tx_done <= 5��    b   '                  �                     5�_�   	              
   c   (    ����                                                                                                                                                                                                                                                                                                                                                             f;x9     �   b   d   �      )                            tx_done <= ''5��    b   (                  �                     5�_�   
                 c   *    ����                                                                                                                                                                                                                                                                                                                                                             f;x:     �   b   d   �      *                            tx_done <= '1'5��    b   *                  �                     5�_�                    g   #    ����                                                                                                                                                                                                                                                                                                                                                             f;x?     �   g   i   �                              �   g   i   �    5��    g                      G                     �    g                     G                    �    g                     `                     �    g                    _                    �    g                    _                    �    g                 	   _             	       5�_�                    h   !    ����                                                                                                                                                                                                                                                                                                                                                             f;xB     �   g   i   �      !                        tx_done <5��    g   !                  h                     5�_�                    h   "    ����                                                                                                                                                                                                                                                                                                                                                             f;xC     �   g   i   �      #                        tx_done <''5��    g   !                  h                     �    g   !                 h                    5�_�                    h   #    ����                                                                                                                                                                                                                                                                                                                                                             f;xD     �   g   i   �      #                        tx_done <= 5��    g   #                  j                     5�_�                    h   $    ����                                                                                                                                                                                                                                                                                                                                                             f;xE     �   g   i   �      %                        tx_done <= ''5��    g   $                  k                     5�_�                    h   &    ����                                                                                                                                                                                                                                                                                                                                                             f;xF     �   g   i   �      &                        tx_done <= '0'5��    g   &                  m                     5�_�                    o   &    ����                                                                                                                                                                                                                                                                                                                                                             f;xI     �   n   o          +                            tx_done <= '1';5��    n                      �      ,               5�_�                    q   &    ����                                                                                                                                                                                                                                                                                                                                                             f;xK     �   p   q          /                                tx_done <= '1';5��    p                      �      0               5�_�                    y   &    ����                                                                                                                                                                                                                                                                                                                                                             f;xN     �   x   y          /                                tx_done <= '0';5��    x                      )      0               5�_�                    J       ����                                                                                                                                                                                                                                                                                                                                                             f;xb     �   I   J          '                        tx_done <= '0';5��    I                      �      (               5�_�                    J        ����                                                                                                                                                                                                                                                                                                                                                             f;xc     �   I   J           5��    I                      �                     5�_�                     W       ����                                                                                                                                                                                                                                                                                                                                                             f;xh    �   V   W          '                        tx_done <= '0';5��    V                      �	      (               5��