Vim�UnDo� ts�N�.~�8"`�&���V���}\Ⱥ+i�   |   	component contador_cm is   $                           fsM    _�                             ����                                                                                                                                                                                                                                                                                                                                                             fs     �                8architecture interface_fd_arch of interface_hcsr04_fd is�                end entity interface_hcsr04_fd;�         |      entity interface_hcsr04_fd is5��                        3                     �                        N                    �       "                 �                    5�_�                     $        ����                                                                                                                                                                                                                                                                                                                                                             fsL    �   [   ]          	medidor: contador_cm�   4   6          	end component contador_cm;�   #   %   |      	component contador_cm is5��    #                    �                    �    4                    #                    �    [   
                 �                    5��