Vim�UnDo� ��Bu���w�qLa����� *\)N]���   \   architecture arch of tb is                             f:j�    _�                        	    ����                                                                                                                                                                                                                                                                                                                                                             f:j�     �         \      entity tb is end;5��       	                  2                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f:j�    �         \      architecture arch of tb is5��                         T                      5��