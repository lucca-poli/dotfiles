Vim�UnDo� �0��+Sr����!t��xh,j�.��(��26   	                                  e�!�    _�                              ����                                                                                                                                                                                                                                                                                                                                                             e�!    �                   �               5��                                                  �                                                �                                                �                                                �                                                �                                                �                                                �                                                �                                                �                                                �                                                �                                                �                                                �                                                �                                              �                                                �                                                �                                                �                                                �                                                �                                                �                                                �                                                  �                                                5��