Vim�UnDo� vg�d.�*(�֭�$z*a&W�{]Y�>�HP�L�   W   >        wait until falling_edge(serial_out) for PERIODOCLK*80;   B   +                       fCn�    _�                        	    ����                                                                                                                                                                                                                                                                                                                                                             f:i�     �         W      entity tb is end;5��       	                  2                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f:i�    �         W      architecture arch of tb is5��                         T                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f:j�     �         W      entity tbb is end;5��                         1                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f:j�    �         W      architecture arch of tbb is5��                         R                      5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                                             fB��     �         W      *    constant PERIODOCLK : time := 20   ns;5��       *                  c                     5�_�                       +    ����                                                                                                                                                                                                                                                                                                                                                             fB��     �         W      0    constant PERIODOCLK : time := 20   ns; 50Mhz5��       +                  d                     5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                                             fB�   	 �         W      *    constant PERIODOBIT : time := 20*4 ns;5��       *                  �                     5�_�                      "    ����                                                                                                                                                                                                                                                                                                                                                             fCaS     �         W      2    constant PERIODOBIT : time := 20*4 ns; -- 5kHz5��       "                  �                     5�_�                      "    ����                                                                                                                                                                                                                                                                                                                                                             fCaY     �         W      0    constant PERIODOBIT : time := *4 ns; -- 5kHz5��       "                 �                    5�_�                       &    ����                                                                                                                                                                                                                                                                                                                                                             fCa]   
 �         W      1    constant PERIODOBIT : time := 0.2 ns; -- 5kHz5��       &                 �                    5�_�                       "    ����                                                                                                                                                                                                                                                                                                                               "          $       v   $    fCdA     �         W      1    constant PERIODOBIT : time := 0.2 ms; -- 5kHz5��       "                 �                    �       $                 �                    5�_�                       &    ����                                                                                                                                                                                                                                                                                                                               "          $       v   $    fCdF     �         W      1    constant PERIODOBIT : time := 208 ms; -- 5kHz5��       &                 �                    5�_�                       .    ����                                                                                                                                                                                                                                                                                                                               "          $       v   $    fCdH     �         W      1    constant PERIODOBIT : time := 208 us; -- 5kHz5��       -                 �                    5�_�                       -    ����                                                                                                                                                                                                                                                                                                                               -          /       v   /    fCe�     �         W      3    constant PERIODOBIT : time := 208 us; -- 4.8kHz5��       -                 �                    5�_�                       $    ����                                                                                                                                                                                                                                                                                                                               -          /       v   /    fCf    �         W      1    constant PERIODOBIT : time := 208 us; -- 5kHz5��       $                 �                    5�_�                     B   +    ����                                                                                                                                                                                                                                                                                                                            B   +       B   <       v   <    fCn�    �   A   C   W      >        wait until falling_edge(serial_out) for PERIODOCLK*80;5��    A   +                  Y
                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             fCaU     �         W          w5��              ,          q      ,              5�_�      	                &    ����                                                                                                                                                                                                                                                                                                                                                             fB�     �         W      1    constant PERIODOBIT : time := 0.2 ns; -- 5kHz5��       "                 �                    5�_�      
           	      &    ����                                                                                                                                                                                                                                                                                                                                                             fB�-    �         W      1    constant PERIODOBIT : time := 0.2 ms; -- 5kHz5��       &                 �                    5�_�   	               
      &    ����                                                                                                                                                                                                                                                                                                                                                             fB�9     �         W      1    constant PERIODOBIT : time := 0.2 us; -- 5kHz5��       &                 �                    5��