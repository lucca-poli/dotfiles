Vim�UnDo� X��f��)��l�����n�R8q�Yp)E                  );            E       E   E   E    f ��    _�                             ����                                                                                                                                                                                                                                                                                                                                                             f �/     �                   �               5��                                          �       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �2     �                e n t i t y multisteps i s5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �2     �                en t i t y multisteps i s5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �3     �                ent i t y multisteps i s5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �3     �                enti t y multisteps i s5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �3     �                entit y multisteps i s5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �7     �                entity multisteps i s5��                                                5�_�      	                      ����                                                                                                                                                                                                                                                                                                                                                             f �:     �               po r t (5��                                                5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                             f �;     �                   po r t (5��                                               5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                             f �<     �                   por t (5��                                               5�_�   
                         ����                                                                                                                                                                                                                                                                                                                                                             f �=     �               clk , r s t : in b i t ;5��                                                 5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �@     �                        clk , r s t : in b i t ;5��                         +                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �A     �                       clk, r s t : in b i t ;5��                         .                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �B     �                       clk, rs t : in b i t ;5��                         /                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �D     �                       clk, rst : in b i t ;5��                         7                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �D     �                       clk, rst : in bi t ;5��                         8                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �E     �                       clk, rst : in bit ;5��                         9                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f �G     �               1msgi : in b i t _ v e c t o r (5 1 1 downto 0 ) ;5��                          ;                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �I     �               9        msgi : in b i t _ v e c t o r (5 1 1 downto 0 ) ;5��                         N                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �I     �               8        msgi : in bi t _ v e c t o r (5 1 1 downto 0 ) ;5��                         O                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �J     �               7        msgi : in bit _ v e c t o r (5 1 1 downto 0 ) ;5��                         P                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �J     �               6        msgi : in bit_ v e c t o r (5 1 1 downto 0 ) ;5��                         Q                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �J     �               5        msgi : in bit_v e c t o r (5 1 1 downto 0 ) ;5��                         R                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �J     �               4        msgi : in bit_ve c t o r (5 1 1 downto 0 ) ;5��                         S                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �J     �               3        msgi : in bit_vec t o r (5 1 1 downto 0 ) ;5��                         T                      5�_�                          ����                                                                                                                                                                                                                                                                                                                                                             f �M     �               2        msgi : in bit_vect o r (5 1 1 downto 0 ) ;5��                         U                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �M     �               1        msgi : in bit_vecto r (5 1 1 downto 0 ) ;5��                         V                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �N     �               0        msgi : in bit_vector (5 1 1 downto 0 ) ;5��                         W                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f �O     �               /        msgi : in bit_vector(5 1 1 downto 0 ) ;5��                         Y                      5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                                             f �O     �               .        msgi : in bit_vector(51 1 downto 0 ) ;5��                         Z                      5�_�       "           !      )    ����                                                                                                                                                                                                                                                                                                                                                             f �R     �               -        msgi : in bit_vector(511 downto 0 ) ;5��       )                  d                      5�_�   !   #           "      *    ����                                                                                                                                                                                                                                                                                                                                                             f �R     �               ,        msgi : in bit_vector(511 downto 0) ;5��       *                  e                      5�_�   "   $           #           ����                                                                                                                                                                                                                                                                                                                                                             f �T     �               2haso : out b i t _ v e c t o r (2 5 5 downto 0 ) ;5��                          g                      5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                                             f �W     �               :        haso : out b i t _ v e c t o r (2 5 5 downto 0 ) ;5��                         {                      5�_�   $   &           %          ����                                                                                                                                                                                                                                                                                                                                                             f �X     �               9        haso : out bi t _ v e c t o r (2 5 5 downto 0 ) ;5��                         |                      5�_�   %   '           &          ����                                                                                                                                                                                                                                                                                                                                                             f �X     �               8        haso : out bit _ v e c t o r (2 5 5 downto 0 ) ;5��                         }                      5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                                             f �X     �               7        haso : out bit_ v e c t o r (2 5 5 downto 0 ) ;5��                         ~                      5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                             f �X     �               6        haso : out bit_v e c t o r (2 5 5 downto 0 ) ;5��                                               5�_�   (   *           )          ����                                                                                                                                                                                                                                                                                                                                                             f �Y     �               5        haso : out bit_ve c t o r (2 5 5 downto 0 ) ;5��                         �                      5�_�   )   +           *          ����                                                                                                                                                                                                                                                                                                                                                             f �Y     �               4        haso : out bit_vec t o r (2 5 5 downto 0 ) ;5��                         �                      5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                                             f �Y     �               3        haso : out bit_vect o r (2 5 5 downto 0 ) ;5��                         �                      5�_�   +   -           ,          ����                                                                                                                                                                                                                                                                                                                                                             f �Y     �               2        haso : out bit_vecto r (2 5 5 downto 0 ) ;5��                         �                      5�_�   ,   .           -          ����                                                                                                                                                                                                                                                                                                                                                             f �Z     �               1        haso : out bit_vector (2 5 5 downto 0 ) ;5��                         �                      5�_�   -   /           .          ����                                                                                                                                                                                                                                                                                                                                                             f �[     �               0        haso : out bit_vector(2 5 5 downto 0 ) ;5��                         �                      5�_�   .   1           /           ����                                                                                                                                                                                                                                                                                                                                                             f �[     �               /        haso : out bit_vector(25 5 downto 0 ) ;5��                          �                      5�_�   /   2   0       1      *    ����                                                                                                                                                                                                                                                                                                                                                             f �a     �               .        haso : out bit_vector(255 downto 0 ) ;5��       *                  �                      5�_�   1   3           2      +    ����                                                                                                                                                                                                                                                                                                                                                             f �c     �               -        haso : out bit_vector(255 downto 0) ;5��       +                  �                      5�_�   2   4           3      +    ����                                                                                                                                                                                                                                                                                                                                                             f �e     �               .        haso : out bit_vector(255 downto 0)l ;5��       +                  �                      5�_�   3   5           4      +    ����                                                                                                                                                                                                                                                                                                                                                             f �e     �               -        haso : out bit_vector(255 downto 0) ;5��       +                  �                      5�_�   4   6           5           ����                                                                                                                                                                                                                                                                                                                                                             f �f     �               done : out b i t5��                          �                      5�_�   5   7           6          ����                                                                                                                                                                                                                                                                                                                                                             f �h     �                       done : out b i t5��                         �                      5�_�   6   8           7          ����                                                                                                                                                                                                                                                                                                                                                             f �i     �                       done : out bi t5��                         �                      5�_�   7   9           8          ����                                                                                                                                                                                                                                                                                                                                                             f �l     �                 ) ;5��                         �                      5�_�   8   :           9           ����                                                                                                                                                                                                                                                                                                                                                             f �m     �                 );5��                          �                      5�_�   9   ;           :          ����                                                                                                                                                                                                                                                                                                                                                             f �o     �                     �               5��                          �                      �                         �                     5�_�   :   <           ;          ����                                                                                                                                                                                                                                                                                                                                                             f ��     �                 end 5��                         �                      �                         �                      �                         �                      �                     
   �              
       �              
          �       
              �                        �                     5�_�   ;   =           <          ����                                                                                                                                                                                                                                                                                                                                                             f ��     �                 end architecture �   	            architecture rtl of  is�                     �   	              arch�                  �               5��                          �                      �                          �                      �    	                      �                      �    	                     �                      �    	                     �                      �    	                     �                      �    	                     �                     �    	                     �                     �    	                     �                     �    	                     �                     �    	                    �                      �                          �                       �                        �                      �                                              �    	                  
   �               
       �                                              5�_�   <   >           =   
       ����                                                                                                                                                                                                                                                                                                                            
          
          v       f ��     �   
          �                 end architecture rtl;�   
          �   
          �   
          �   
          �   
          �   
          �   
          �   
          �   
          �   
          �   
          �   	            !architecture rtl of multisteps is5��    	                    �                     �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                     	                	       �    	                     �                      �              	       
         	       
       5�_�   =   ?           >          ����                                                                                                                                                                                                                                                                                                                            
   $       
          v       f ��     �   
                �   
          5��    
                      �                      �    
                      �                      �    
                     �                      �                      
   �               
       5�_�   >   @           ?           ����                                                                                                                                                                                                                                                                                                                                                V       f ��     �             �             �                    component 5��                          �                      �                          �               �       5�_�   ?   A           @          ����                                                                                                                                                                                                                                                                                                                                                 V       f ��     �                   component ch is5��                         �                      5�_�   @   B           A          ����                                                                                                                                                                                                                                                                                                                                                 V       f ��     �                   component  is�             5��                         �                      5�_�   A   C           B          ����                                                                                                                                                                                                                                                                                                                                               V       f ��     �               0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)5��       0                F                    5�_�   B   D           C          ����                                                                                                                                                                                                                                                                                                                             	                 V       f ��     �             �             �                        port (   O            x, y, z: in bit_vector(31 downto 0); q: out bit_vector(31 downto 0)   
        );5��                                j               �                                        �       5�_�   C   E           D          ����                                                                                                                                                                                                                                                                                                                                                      f ��     �               @    	ai, bi, ci, di, ei, fi, gi, hi: in bit_vector(31 downto 0);   (        kpw: in bit_vector(31 downto 0);   C        ao, bo, co, do, eo, fo, go, ho: out bit_vector(31 downto 0)   
        );�               
    port (5��                                              �                                              �                         _                     �                         �                     �                         �                     5�_�   D               E          ����                                                                                                                                                                                                                                                                                                                                                      f ��    �                           );5��                         �                     5�_�   /           1   0      !    ����                                                                                                                                                                                                                                                                                                                                                             f �\     �               -        haso : out bit_vector(255downto 0 ) ;5��       !                  �                      5�_�                          ����                                                                                                                                                                                                                                                                                                                                                             f �K     �               1        msgi : in bit_vect  r (5 1 1 downto 0 ) ;5��                         V                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f �K     �               0        msgi : in bit_vect   (5 1 1 downto 0 ) ;5��                         W                      5��