Vim�UnDo� ��]ia=,�:�XQg���4�r�����:�)JK   V   L            assert false report integer'image(HEXA*iteration) severity note;   P   .                   f�   4 _�                             ����                                                                                                                                                                                                                                                                                                                                                             f �/     �                   �               5��                                          �       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �2     �                e n t i t y multisteps i s5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �2     �                en t i t y multisteps i s5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �3     �                ent i t y multisteps i s5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �3     �                enti t y multisteps i s5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �3     �                entit y multisteps i s5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �7     �                entity multisteps i s5��                                                5�_�      	                      ����                                                                                                                                                                                                                                                                                                                                                             f �:     �               po r t (5��                                                5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                             f �;     �                   po r t (5��                                               5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                             f �<     �                   por t (5��                                               5�_�   
                         ����                                                                                                                                                                                                                                                                                                                                                             f �=     �               clk , r s t : in b i t ;5��                                                 5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �@     �                        clk , r s t : in b i t ;5��                         +                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �A     �                       clk, r s t : in b i t ;5��                         .                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �B     �                       clk, rs t : in b i t ;5��                         /                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �D     �                       clk, rst : in b i t ;5��                         7                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �D     �                       clk, rst : in bi t ;5��                         8                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �E     �                       clk, rst : in bit ;5��                         9                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f �G     �               1msgi : in b i t _ v e c t o r (5 1 1 downto 0 ) ;5��                          ;                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �I     �               9        msgi : in b i t _ v e c t o r (5 1 1 downto 0 ) ;5��                         N                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �I     �               8        msgi : in bi t _ v e c t o r (5 1 1 downto 0 ) ;5��                         O                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �J     �               7        msgi : in bit _ v e c t o r (5 1 1 downto 0 ) ;5��                         P                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �J     �               6        msgi : in bit_ v e c t o r (5 1 1 downto 0 ) ;5��                         Q                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �J     �               5        msgi : in bit_v e c t o r (5 1 1 downto 0 ) ;5��                         R                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �J     �               4        msgi : in bit_ve c t o r (5 1 1 downto 0 ) ;5��                         S                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �J     �               3        msgi : in bit_vec t o r (5 1 1 downto 0 ) ;5��                         T                      5�_�                          ����                                                                                                                                                                                                                                                                                                                                                             f �M     �               2        msgi : in bit_vect o r (5 1 1 downto 0 ) ;5��                         U                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �M     �               1        msgi : in bit_vecto r (5 1 1 downto 0 ) ;5��                         V                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f �N     �               0        msgi : in bit_vector (5 1 1 downto 0 ) ;5��                         W                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f �O     �               /        msgi : in bit_vector(5 1 1 downto 0 ) ;5��                         Y                      5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                                             f �O     �               .        msgi : in bit_vector(51 1 downto 0 ) ;5��                         Z                      5�_�       "           !      )    ����                                                                                                                                                                                                                                                                                                                                                             f �R     �               -        msgi : in bit_vector(511 downto 0 ) ;5��       )                  d                      5�_�   !   #           "      *    ����                                                                                                                                                                                                                                                                                                                                                             f �R     �               ,        msgi : in bit_vector(511 downto 0) ;5��       *                  e                      5�_�   "   $           #           ����                                                                                                                                                                                                                                                                                                                                                             f �T     �               2haso : out b i t _ v e c t o r (2 5 5 downto 0 ) ;5��                          g                      5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                                             f �W     �               :        haso : out b i t _ v e c t o r (2 5 5 downto 0 ) ;5��                         {                      5�_�   $   &           %          ����                                                                                                                                                                                                                                                                                                                                                             f �X     �               9        haso : out bi t _ v e c t o r (2 5 5 downto 0 ) ;5��                         |                      5�_�   %   '           &          ����                                                                                                                                                                                                                                                                                                                                                             f �X     �               8        haso : out bit _ v e c t o r (2 5 5 downto 0 ) ;5��                         }                      5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                                             f �X     �               7        haso : out bit_ v e c t o r (2 5 5 downto 0 ) ;5��                         ~                      5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                             f �X     �               6        haso : out bit_v e c t o r (2 5 5 downto 0 ) ;5��                                               5�_�   (   *           )          ����                                                                                                                                                                                                                                                                                                                                                             f �Y     �               5        haso : out bit_ve c t o r (2 5 5 downto 0 ) ;5��                         �                      5�_�   )   +           *          ����                                                                                                                                                                                                                                                                                                                                                             f �Y     �               4        haso : out bit_vec t o r (2 5 5 downto 0 ) ;5��                         �                      5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                                             f �Y     �               3        haso : out bit_vect o r (2 5 5 downto 0 ) ;5��                         �                      5�_�   +   -           ,          ����                                                                                                                                                                                                                                                                                                                                                             f �Y     �               2        haso : out bit_vecto r (2 5 5 downto 0 ) ;5��                         �                      5�_�   ,   .           -          ����                                                                                                                                                                                                                                                                                                                                                             f �Z     �               1        haso : out bit_vector (2 5 5 downto 0 ) ;5��                         �                      5�_�   -   /           .          ����                                                                                                                                                                                                                                                                                                                                                             f �[     �               0        haso : out bit_vector(2 5 5 downto 0 ) ;5��                         �                      5�_�   .   1           /           ����                                                                                                                                                                                                                                                                                                                                                             f �[     �               /        haso : out bit_vector(25 5 downto 0 ) ;5��                          �                      5�_�   /   2   0       1      *    ����                                                                                                                                                                                                                                                                                                                                                             f �a     �               .        haso : out bit_vector(255 downto 0 ) ;5��       *                  �                      5�_�   1   3           2      +    ����                                                                                                                                                                                                                                                                                                                                                             f �c     �               -        haso : out bit_vector(255 downto 0) ;5��       +                  �                      5�_�   2   4           3      +    ����                                                                                                                                                                                                                                                                                                                                                             f �e     �               .        haso : out bit_vector(255 downto 0)l ;5��       +                  �                      5�_�   3   5           4      +    ����                                                                                                                                                                                                                                                                                                                                                             f �e     �               -        haso : out bit_vector(255 downto 0) ;5��       +                  �                      5�_�   4   6           5           ����                                                                                                                                                                                                                                                                                                                                                             f �f     �               done : out b i t5��                          �                      5�_�   5   7           6          ����                                                                                                                                                                                                                                                                                                                                                             f �h     �                       done : out b i t5��                         �                      5�_�   6   8           7          ����                                                                                                                                                                                                                                                                                                                                                             f �i     �                       done : out bi t5��                         �                      5�_�   7   9           8          ����                                                                                                                                                                                                                                                                                                                                                             f �l     �                 ) ;5��                         �                      5�_�   8   :           9           ����                                                                                                                                                                                                                                                                                                                                                             f �m     �                 );5��                          �                      5�_�   9   ;           :          ����                                                                                                                                                                                                                                                                                                                                                             f �o     �                     �               5��                          �                      �                         �                     5�_�   :   <           ;          ����                                                                                                                                                                                                                                                                                                                                                             f ��     �                 end 5��                         �                      �                         �                      �                         �                      �                     
   �              
       �              
          �       
              �                        �                     5�_�   ;   =           <          ����                                                                                                                                                                                                                                                                                                                                                             f ��     �                 end architecture �   	            architecture rtl of  is�                     �   	              arch�                  �               5��                          �                      �                          �                      �    	                      �                      �    	                     �                      �    	                     �                      �    	                     �                      �    	                     �                     �    	                     �                     �    	                     �                     �    	                     �                     �    	                    �                      �                          �                       �                        �                      �                                              �    	                  
   �               
       �                                              5�_�   <   >           =   
       ����                                                                                                                                                                                                                                                                                                                            
          
          v       f ��     �   
          �                 end architecture rtl;�   
          �   
          �   
          �   
          �   
          �   
          �   
          �   
          �   
          �   
          �   
          �   	            !architecture rtl of multisteps is5��    	                    �                     �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                                            �    	                     �                      �                     	                	       �    	                     �                      �              	       
         	       
       5�_�   =   ?           >          ����                                                                                                                                                                                                                                                                                                                            
   $       
          v       f ��     �   
                �   
          5��    
                      �                      �    
                      �                      �    
                     �                      �                      
   �               
       5�_�   >   @           ?           ����                                                                                                                                                                                                                                                                                                                                                V       f ��     �             �             �                    component 5��                          �                      �                          �               �       5�_�   ?   A           @          ����                                                                                                                                                                                                                                                                                                                                                 V       f ��     �                   component ch is5��                         �                      5�_�   @   B           A          ����                                                                                                                                                                                                                                                                                                                                                 V       f ��     �                   component  is�             5��                         �                      5�_�   A   C           B          ����                                                                                                                                                                                                                                                                                                                                               V       f ��     �               0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)5��       0                F                    5�_�   B   D           C          ����                                                                                                                                                                                                                                                                                                                             	                 V       f ��     �             �             �                        port (   O            x, y, z: in bit_vector(31 downto 0); q: out bit_vector(31 downto 0)   
        );5��                                j               �                                        �       5�_�   C   E           D          ����                                                                                                                                                                                                                                                                                                                                                      f ��     �               @    	ai, bi, ci, di, ei, fi, gi, hi: in bit_vector(31 downto 0);   (        kpw: in bit_vector(31 downto 0);   C        ao, bo, co, do, eo, fo, go, ho: out bit_vector(31 downto 0)   
        );�               
    port (5��                                              �                                              �                         _                     �                         �                     �                         �                     5�_�   D   F           E          ����                                                                                                                                                                                                                                                                                                                                                      f ��    �                           );5��                         �                     5�_�   E   G           F           ����                                                                                                                                                                                                                                                                                                                                                      f ��     �                   �             5��                          �                     �                          �                     �                         �                     �                         �                     5�_�   F   H           G          ����                                                                                                                                                                                                                                                                                                                                                      f ��     �                   �             �             5��                                                �                                      �       5�_�   G   I           H      	    ����                                                                                                                                                                                                                                                                                                                                                      f ��     �               !    type constants_type is record5��       	                 	                    5�_�   H   J           I          ����                                                                                                                                                                                                                                                                                                                                                      f ��     �                       CONSTANT_1 : integer;5��              
          $      
              5�_�   I   L           J          ����                                                                                                                                                                                                                                                                                                                                                      f ��     �                        CONSTANT_2 : integer;5��                          3                     5�_�   J   N   K       L          ����                                                                                                                                                                                                                                                                                                                                                      f ��     �      V       �             5��                   ?       3              �      5�_�   L   O   M       N      
    ����                                                                                                                                                                                                                                                                                                                              
       U   
          
    f �D     �      V   ]   ?           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;           H_0 : integer;5��       
                 =                    �       
                 T                    �       
                 k                    �       
                 �                    �       
                 �                    �       
                 �                    �       
                 �                    �       
                 �                    �       
                 �                    �       
                                     �        
                 $                    �    !   
                 <                    �    "   
                 T                    �    #   
                 l                    �    $   
                 �                    �    %   
                 �                    �    &   
                 �                    �    '   
                 �                    �    (   
                 �                    �    )   
                 �                    �    *   
                                     �    +   
                 ,                    �    ,   
                 D                    �    -   
                 \                    �    .   
                 t                    �    /   
                 �                    �    0   
                 �                    �    1   
                 �                    �    2   
                 �                    �    3   
                 �                    �    4   
                                     �    5   
                                     �    6   
                 4                    �    7   
                 L                    �    8   
                 d                    �    9   
                 |                    �    :   
                 �                    �    ;   
                 �                    �    <   
                 �                    �    =   
                 �                    �    >   
                 �                    �    ?   
                                     �    @   
                 $                    �    A   
                 <                    �    B   
                 T                    �    C   
                 l                    �    D   
                 �                    �    E   
                 �                    �    F   
                 �                    �    G   
                 �                    �    H   
                 �                    �    I   
                 �                    �    J   
                                     �    K   
                 ,                    �    L   
                 D                    �    M   
                 \                    �    N   
                 t                    �    O   
                 �                    �    P   
                 �                    �    Q   
                 �                    �    R   
                 �                    �    S   
                 �                    �    T   
                                     5�_�   N   P           O   V   
    ����                                                                                                                                                                                                                                                                                                                              
       U   
          
    f �J     �   U   V          *        -- Define more constants as needed5��    U                            +               5�_�   O   Q           P   W       ����                                                                                                                                                                                                                                                                                                                           V   
          
       V   
    f �Z     �   W   Y   \    5��    W                      '                     �    W                      '                     5�_�   P   R           Q   W       ����                                                                                                                                                                                                                                                                                                                           V   
          
       V   
    f �[     �   W   �   ]    �   W   X   ]    5��    W               B       '              "      5�_�   Q   S           R   X   	    ����                                                                                                                                                                                                                                                                                                                           V   
          
       V   
    f �l     �   W   Y   �          type h_vector is record5��    W   	                 0                    5�_�   R   T           S   X   	    ����                                                                                                                                                                                                                                                                                                                           V   
          
       V   
    f ��     �   W   Y   �          type k_vector is record5��    W   	                 0                    5�_�   S   U           T   a        ����                                                                                                                                                                                                                                                                                                                           a   	       �   	       V   	    f ��     �   `   a       8           H_8 : integer;           H_9 : integer;           H_10 : integer;           H_11 : integer;           H_12 : integer;           H_13 : integer;           H_14 : integer;           H_15 : integer;           H_16 : integer;           H_17 : integer;           H_18 : integer;           H_19 : integer;           H_20 : integer;           H_21 : integer;           H_22 : integer;           H_23 : integer;           H_24 : integer;           H_25 : integer;           H_26 : integer;           H_27 : integer;           H_28 : integer;           H_29 : integer;           H_30 : integer;           H_31 : integer;           H_32 : integer;           H_33 : integer;           H_34 : integer;           H_35 : integer;           H_36 : integer;           H_37 : integer;           H_38 : integer;           H_39 : integer;           H_40 : integer;           H_41 : integer;           H_42 : integer;           H_43 : integer;           H_44 : integer;           H_45 : integer;           H_46 : integer;           H_47 : integer;           H_48 : integer;           H_49 : integer;           H_50 : integer;           H_51 : integer;           H_52 : integer;           H_53 : integer;           H_54 : integer;           H_55 : integer;           H_56 : integer;           H_57 : integer;           H_58 : integer;           H_59 : integer;           H_60 : integer;           H_61 : integer;           H_62 : integer;           H_63 : integer;5��    `       8               �      >              5�_�   T   V           U           ����                                                                                                                                                                                                                                                                                                                           U   	          	       V   	    f ��     �   T   V                  H_63 : integer;�   S   U                  H_62 : integer;�   R   T                  H_61 : integer;�   Q   S                  H_60 : integer;�   P   R                  H_59 : integer;�   O   Q                  H_58 : integer;�   N   P                  H_57 : integer;�   M   O                  H_56 : integer;�   L   N                  H_55 : integer;�   K   M                  H_54 : integer;�   J   L                  H_53 : integer;�   I   K                  H_52 : integer;�   H   J                  H_51 : integer;�   G   I                  H_50 : integer;�   F   H                  H_49 : integer;�   E   G                  H_48 : integer;�   D   F                  H_47 : integer;�   C   E                  H_46 : integer;�   B   D                  H_45 : integer;�   A   C                  H_44 : integer;�   @   B                  H_43 : integer;�   ?   A                  H_42 : integer;�   >   @                  H_41 : integer;�   =   ?                  H_40 : integer;�   <   >                  H_39 : integer;�   ;   =                  H_38 : integer;�   :   <                  H_37 : integer;�   9   ;                  H_36 : integer;�   8   :                  H_35 : integer;�   7   9                  H_34 : integer;�   6   8                  H_33 : integer;�   5   7                  H_32 : integer;�   4   6                  H_31 : integer;�   3   5                  H_30 : integer;�   2   4                  H_29 : integer;�   1   3                  H_28 : integer;�   0   2                  H_27 : integer;�   /   1                  H_26 : integer;�   .   0                  H_25 : integer;�   -   /                  H_24 : integer;�   ,   .                  H_23 : integer;�   +   -                  H_22 : integer;�   *   ,                  H_21 : integer;�   )   +                  H_20 : integer;�   (   *                  H_19 : integer;�   '   )                  H_18 : integer;�   &   (                  H_17 : integer;�   %   '                  H_16 : integer;�   $   &                  H_15 : integer;�   #   %                  H_14 : integer;�   "   $                  H_13 : integer;�   !   #                  H_12 : integer;�       "                  H_11 : integer;�      !                  H_10 : integer;�                         H_9 : integer;�                        H_8 : integer;�                        H_7 : integer;�                        H_6 : integer;�                        H_5 : integer;�                        H_4 : integer;�                        H_3 : integer;�                        H_2 : integer;�                        H_1 : integer;�         g              H_0 : integer;5��                        $                    �                        ;                    �                        R                    �                        i                    �                        �                    �                        �                    �                        �                    �                        �                    �                        �                    �                        �                    �                        
                    �                         "                    �    !                    :                    �    "                    R                    �    #                    j                    �    $                    �                    �    %                    �                    �    &                    �                    �    '                    �                    �    (                    �                    �    )                    �                    �    *                                        �    +                    *                    �    ,                    B                    �    -                    Z                    �    .                    r                    �    /                    �                    �    0                    �                    �    1                    �                    �    2                    �                    �    3                    �                    �    4                                        �    5                                        �    6                    2                    �    7                    J                    �    8                    b                    �    9                    z                    �    :                    �                    �    ;                    �                    �    <                    �                    �    =                    �                    �    >                    �                    �    ?                    
                    �    @                    "                    �    A                    :                    �    B                    R                    �    C                    j                    �    D                    �                    �    E                    �                    �    F                    �                    �    G                    �                    �    H                    �                    �    I                    �                    �    J                                        �    K                    *                    �    L                    B                    �    M                    Z                    �    N                    r                    �    O                    �                    �    P                    �                    �    Q                    �                    �    R                    �                    �    S                    �                    �    T                                        5�_�   U   Y           V      	    ����                                                                                                                                                                                                                                                                                                                           U   	          	       V   	    f ��     �         g          type h_vector is record5��       	                 	                    5�_�   V   Z   X       Y           ����                                                                                                                                                                                                                                                                                                                                      a           V        f ��     �   _   a                  H_7 : integer;�   ^   `                  H_6 : integer;�   ]   _                  H_5 : integer;�   \   ^                  H_4 : integer;�   [   ]                  H_3 : integer;�   Z   \                  H_2 : integer;�   Y   [                  H_1 : integer;�   X   Z                  H_0 : integer;�   T   V                  K_63 : integer;�   S   U                  K_62 : integer;�   R   T                  K_61 : integer;�   Q   S                  K_60 : integer;�   P   R                  K_59 : integer;�   O   Q                  K_58 : integer;�   N   P                  K_57 : integer;�   M   O                  K_56 : integer;�   L   N                  K_55 : integer;�   K   M                  K_54 : integer;�   J   L                  K_53 : integer;�   I   K                  K_52 : integer;�   H   J                  K_51 : integer;�   G   I                  K_50 : integer;�   F   H                  K_49 : integer;�   E   G                  K_48 : integer;�   D   F                  K_47 : integer;�   C   E                  K_46 : integer;�   B   D                  K_45 : integer;�   A   C                  K_44 : integer;�   @   B                  K_43 : integer;�   ?   A                  K_42 : integer;�   >   @                  K_41 : integer;�   =   ?                  K_40 : integer;�   <   >                  K_39 : integer;�   ;   =                  K_38 : integer;�   :   <                  K_37 : integer;�   9   ;                  K_36 : integer;�   8   :                  K_35 : integer;�   7   9                  K_34 : integer;�   6   8                  K_33 : integer;�   5   7                  K_32 : integer;�   4   6                  K_31 : integer;�   3   5                  K_30 : integer;�   2   4                  K_29 : integer;�   1   3                  K_28 : integer;�   0   2                  K_27 : integer;�   /   1                  K_26 : integer;�   .   0                  K_25 : integer;�   -   /                  K_24 : integer;�   ,   .                  K_23 : integer;�   +   -                  K_22 : integer;�   *   ,                  K_21 : integer;�   )   +                  K_20 : integer;�   (   *                  K_19 : integer;�   '   )                  K_18 : integer;�   &   (                  K_17 : integer;�   %   '                  K_16 : integer;�   $   &                  K_15 : integer;�   #   %                  K_14 : integer;�   "   $                  K_13 : integer;�   !   #                  K_12 : integer;�       "                  K_11 : integer;�      !                  K_10 : integer;�                         K_9 : integer;�                        K_8 : integer;�                        K_7 : integer;�                        K_6 : integer;�                        K_5 : integer;�                        K_4 : integer;�                        K_3 : integer;�                        K_2 : integer;�                        K_1 : integer;�         g              K_0 : integer;5��                        *                    �                        Q                    �                        x                    �                        �                    �                        �                    �                        �                    �                                            �                        ;                    �                        b                    �                        �                    �                        �                    �                         �                    �    !                                        �    "                    )                    �    #                    Q                    �    $                    y                    �    %                    �                    �    &                    �                    �    '                    �                    �    (                                        �    )                    A                    �    *                    i                    �    +                    �                    �    ,                    �                    �    -                    �                    �    .                    	                    �    /                    1                    �    0                    Y                    �    1                    �                    �    2                    �                    �    3                    �                    �    4                    �                    �    5                    !                    �    6                    I                    �    7                    q                    �    8                    �                    �    9                    �                    �    :                    �                    �    ;                                        �    <                    9                    �    =                    a                    �    >                    �                    �    ?                    �                    �    @                    �                    �    A                    	                    �    B                    )	                    �    C                    Q	                    �    D                    y	                    �    E                    �	                    �    F                    �	                    �    G                    �	                    �    H                    
                    �    I                    A
                    �    J                    i
                    �    K                    �
                    �    L                    �
                    �    M                    �
                    �    N                    	                    �    O                    1                    �    P                    Y                    �    Q                    �                    �    R                    �                    �    S                    �                    �    T                    �                    �    X                    Q                    �    Y                    x                    �    Z                    �                    �    [                    �                    �    \                    �                    �    ]                                        �    ^                    ;                    �    _                    b                    5�_�   Y   \           Z   a       ����                                                                                                                                                                                                                                                                                                                                      a           V        f �     �   a   c   g    5��    a                      �                     �    a                      �                     5�_�   Z   ]   [       \   b        ����                                                                                                                                                                                                                                                                                                                                      a           V        f �     �   b   h   i          �   c   d   i    �   b   d   h    5��    b                      �                     �    b                      �                     �    b                    �              �       5�_�   \   ^           ]   c       ����                                                                                                                                                                                                                                                                                                                                      a           V        f �     �   b   d   m      ,    constant CONSTANTS : constants_type := (5��    b          	          �      	              5�_�   ]   _           ^   c       ����                                                                                                                                                                                                                                                                                                                                      a           V        f �      �   b   d   m      $    constant H : constants_type := (5��    b                    �                    �    b                    �                    �    b                    �                    �    b                    �                    5�_�   ^   `           _   c        ����                                                                                                                                                                                                                                                                                                                           Y          `          V       f �-     �   c   l   m    �   c   d   m    5��    c                      �              8      5�_�   _   a           `   d        ����                                                                                                                                                                                                                                                                                                                           d          k          V       f �>     �   j   l          &        H_7 : bit_vector(31 downto 0);�   i   k          &        H_6 : bit_vector(31 downto 0);�   h   j          &        H_5 : bit_vector(31 downto 0);�   g   i          &        H_4 : bit_vector(31 downto 0);�   f   h          &        H_3 : bit_vector(31 downto 0);�   e   g          &        H_2 : bit_vector(31 downto 0);�   d   f          &        H_1 : bit_vector(31 downto 0);�   c   e   u      &        H_0 : bit_vector(31 downto 0);5��    c                    �                    �    d                    �                    �    e                                        �    f                    /                    �    g                    W                    �    h                                        �    i                    �                    �    j                    �                    5�_�   `   b           a   d        ����                                                                                                                                                                                                                                                                                                                           k          d          V       f ��     �   j   l          '        H_7 => bit_vector(31 downto 0);�   i   k          '        H_6 => bit_vector(31 downto 0);�   h   j          '        H_5 => bit_vector(31 downto 0);�   g   i          '        H_4 => bit_vector(31 downto 0);�   f   h          '        H_3 => bit_vector(31 downto 0);�   e   g          '        H_2 => bit_vector(31 downto 0);�   d   f          '        H_1 => bit_vector(31 downto 0);�   c   e   u      '        H_0 => bit_vector(31 downto 0);5��    c                    �                    �    d                    �                    �    e                    �                    �    f                    �                    �    g                    �                    �    h                                        �    i                                         �    j                    1                    5�_�   a   c           b   l       ����                                                                                                                                                                                                                                                                                                                           k          d          V       f ��     �   k   l                  CONSTANT_1 => 42,           CONSTANT_2 => 100,5��    k                      3      5               5�_�   b   d           c   l       ����                                                                                                                                                                                                                                                                                                                           k          d          V       f ��     �   k   l          .        -- Initialize more constants as needed5��    k                      3      /               5�_�   c   e           d   d       ����                                                                                                                                                                                                                                                                                                                           k          d          V       f ��     �   c   e   s          �   d   e   s    �   c   e   r    5��    c                      �              	       �    c                  K   �             K       5�_�   d   f           e   d       ����                                                                                                                                                                                                                                                                                                                           l          e          V       f �     �   c   e   s      K    6a09e667 bb67ae85 3c6ef372 a54ff53a 510e527f 9b05688c 1f83d9ab 5be0cd195��    c          G           �      G               5�_�   e   g           f   e       ����                                                                                                                                                                                                                                                                                                                           l          e          V       f �     �   d   f   s              H_0 => ,�   e   f   s    5��    d                  G   �              G       5�_�   f   k           g   d       ����                                                                                                                                                                                                                                                                                                                           l          e          V       f �	     �   c   d              5��    c                      �                     5�_�   g   l   h       k   d       ����                                                                                                                                                                                                                                                                                                                           k          d          V       f �_     �   c   e   r      W        H_0 => 6a09e667 bb67ae85 3c6ef372 a54ff53a 510e527f 9b05688c 1f83d9ab 5be0cd19,5��    c                     �                     5�_�   k   m           l   d       ����                                                                                                                                                                                                                                                                                                                           k          d          V       f �a     �   c   e   r      V        H_0 => 6a09e667bb67ae85 3c6ef372 a54ff53a 510e527f 9b05688c 1f83d9ab 5be0cd19,5��    c          >           �      >               5�_�   l   n           m   e       ����                                                                                                                                                                                                                                                                                                                           k          d          V       f �h     �   d   f   r              H_1 => ,�   e   f   r    5��    d                  >   �              >       5�_�   m   o           n   e       ����                                                                                                                                                                                                                                                                                                                           k          d          V       f �k     �   e   g   r              H_2 => ,�   f   g   r    �   d   f   r      N        H_1 => bb67ae85 3c6ef372 a54ff53a 510e527f 9b05688c 1f83d9ab 5be0cd19,5��    d                     �                     �    d          5           �      5               �    e                  5   �              5       5�_�   n   p           o   f       ����                                                                                                                                                                                                                                                                                                                           k          d          V       f �s     �   j   l   r              H_7 => ,�   k   l   r    �   i   k   r              H_6 => ,�   j   k   r    �   h   j   r              H_5 => ,�   i   j   r    �   g   i   r              H_4 => ,�   h   i   r    �   f   h   r              H_3 => ,�   g   h   r    �   e   g   r      E        H_2 => 3c6ef372 a54ff53a 510e527f 9b05688c 1f83d9ab 5be0cd19,5��    e                     �                     �    e          ,           �      ,               �    f                  ,                 ,       �    f          $                 $               �    g                  #                 #       �    g                     &                     �    h                     7                     �    h                     ?                     �    i                     P                     �    i          	           X      	               �    j                     i                     5�_�   o   q           p   d       ����                                                                                                                                                                                                                                                                                                                           d          k                 f ��     �   d   l   r              H_1 => bb67ae85,           H_2 => 3c6ef372,           H_3 => a54ff53a,           H_4 => 510e527f,           H_5 => 9b05688c,           H_6 => 1f83d9ab,           H_7 => 5be0cd19,�   c   e   r              H_0 => 6a09e667,5��    c                     �                     �    d                     �                     �    e                     �                     �    f                                          �    g                     *                     �    h                     F                     �    i                     b                     �    j                     ~                     5�_�   p   s           q   d       ����                                                                                                                                                                                                                                                                                                                           d          k                 f ��     �   d   l   r              H_1 => 16#bb67ae85,           H_2 => 16#3c6ef372,           H_3 => 16#a54ff53a,           H_4 => 16#510e527f,           H_5 => 16#9b05688c,           H_6 => 16#1f83d9ab,           H_7 => 16#5be0cd19,�   c   e   r              H_0 => 16#6a09e667,5��    c                     �                     �    d                     �                     �    e                     �                     �    f                                          �    g                     9                     �    h                     V                     �    i                     s                     �    j                     �                     5�_�   q   t   r       s   d       ����                                                                                                                                                                                                                                                                                                                           d          k                 f ��     �   c   e   r              H_0 => 16#6a09e667#,5��    c                     �                     5�_�   s   u           t   d       ����                                                                                                                                                                                                                                                                                                                           d          k                 f ��     �   c   e   r              H_0 => (16#6a09e667#,5��    c                     �                    5�_�   t   v           u   d       ����                                                                                                                                                                                                                                                                                                                           d          k                 f ��     �   c   e   r              H_0 => (16#6a09e667#),5��    c                     �                     �    c                 	   �             	       5�_�   u   w           v   d       ����                                                                                                                                                                                                                                                                                                                           d          k                 f ��     �   c   e   r      )        H_0 => to_unsigned(16#6a09e667#),5��    c                    �                    �    c                    �                    5�_�   v   x           w   k       ����                                                                                                                                                                                                                                                                                                                           d          k                 f ��     �   j   l   r              H_7 => 16#5be0cd19#,5��    j                     �                     5�_�   w   y           x          ����                                                                                                                                                                                                                                                                                                                           d          k                 f �     �          s       �         s    �          r    5��                                                  �                                          D       5�_�   x   z           y          ����                                                                                                                                                                                                                                                                                                                           g          n                 f �     �         u    5��                          E                      5�_�   y   {           z      	    ����                                                                                                                                                                                                                                                                                                                           h          o                 f �!     �         v      use IEEE.NUMERIC_STD.ALL;5��       	                 4                     �                         6                      �       
                  5                      �       	                 4                     �       	                 4                     �       	                 4                     �       	                 4                     �       	                 4                     �       	                 4                     �       	                 4                     �       	                 4                     �       	                 4                     �       	                 4                     5�_�   z   |           {   h       ����                                                                                                                                                                                                                                                                                                                           h          o                 f �Y     �   g   i   v      *        H_0 => to_bitvector(16#6a09e667#),5��    g                                           5�_�   {   }           |   h       ����                                                                                                                                                                                                                                                                                                                           h          o                 f �Y     �   g   i   v      )        H_0 => o_bitvector(16#6a09e667#),5��    g                                           5�_�   |   ~           }   h       ����                                                                                                                                                                                                                                                                                                                           h          o                 f �Z     �   g   i   v      (        H_0 => _bitvector(16#6a09e667#),5��    g                                           5�_�   }              ~   h       ����                                                                                                                                                                                                                                                                                                                           h          o                 f �[     �   g   i   v      '        H_0 => bitvector(16#6a09e667#),�   h   i   v    5��    g                                          5�_�   ~   �              h       ����                                                                                                                                                                                                                                                                                                                           h          o                 f �d     �   g   i   v      (        H_0 => bit_vector(16#6a09e667#),5��    g                                          �    g   $                                     5�_�      �           �   h   &    ����                                                                                                                                                                                                                                                                                                                           h          o                 f �l     �   g   i   v      4        H_0 => bit_vector(to_unsigned(16#6a09e667#),5��    g                     �      5       6       5�_�   �   �           �   h       ����                                                                                                                                                                                                                                                                                                                           h          o                 f ��     �   g   i   v      5        H_0 => bit_vector(to_unsigned(16#6a09e667#)),5��    g                                          5�_�   �   �           �   h       ����                                                                                                                                                                                                                                                                                                                           h          o                 f ��     �   g   i   v      4        H_0 => bit_vector(o_unsigned(16#6a09e667#)),5��    g                                          5�_�   �   �           �   h       ����                                                                                                                                                                                                                                                                                                                           h          o                 f ��     �   g   i   v      3        H_0 => bit_vector(_unsigned(16#6a09e667#)),5��    g                                          5�_�   �   �   �       �   v       ����                                                                                                                                                                                                                                                                                                                           h          o                 f ��     �   w               �   x            �   v               �   v            5��    v                      (                     �    v                      (                     �    w               	      )              E      5�_�   �   �           �   w        ����                                                                                                                                                                                                                                                                                                                                               V       f ��     �   w   {   �    �   w   x   �    5��    w                      )              E       5�_�   �   �           �   z        ����                                                                                                                                                                                                                                                                                                                                               V       f ��     �   z   |   �    5��    z                      n                     5�_�   �   �           �   x        ����                                                                                                                                                                                                                                                                                                                           |           �           V        f �     �   w   x          library IEEE;   use IEEE.STD_LOGIC_1164.ALL;   use IEEE.NUMERIC_BIT.ALL;    5��    w                      )      F               5�_�   �   �           �   x        ����                                                                                                                                                                                                                                                                                                                           x           �           V        f �     �   w   x       
   Tfunction convert_to_bit_vector(size : natural; value : integer) return bit_vector is   G    variable result : bit_vector(size - 1 downto 0) := (others => '0');   begin       for i in 0 to size - 1 loop   %        if value and (2**i) /= 0 then               result(i) := '1';           end if;       end loop;       return result;   end function;5��    w       
               )      F              5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                           x           x           V        f �!     �         w    �         w    5��                   
       2              F      5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                #           �           �           V        f �"     �         �    5��                          2                     �                          2                     �                          2                     5�_�   �   �           �      	    ����                                                                                                                                                                                                                                                                                                                $              	                 v       f �&     �         �      Tfunction convert_to_bit_vector(size : natural; value : integer) return bit_vector is5��       	                  <                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                $              	                 v       f �)     �         �      Lfunction to_bit_vector(size : natural; value : integer) return bit_vector is5��                         B                     5�_�   �   �   �       �          ����                                                                                                                                                                                                                                                                                                                $              	                 v       f �Q     �         �      %        if value and (2**i) /= 0 then5��                                              5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                $              	                 v       f �T     �         �      '        if value and ()(2**i) /= 0 then5��                         �      (       (       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f ��     �         �      '        if value and ((2**i) /= 0) then�         �    5��                        �                    5�_�   �   �           �   s       ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f �I     �   r   t   �      2        H_0 => bit_vector(unsigned(16#6a09e667#)),5��    r                     @                     5�_�   �   �           �   s       ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f �K     �   r   t   �      5        H_0 => to_bit_vector(unsigned(16#6a09e667#)),5��    r                     F                     5�_�   �   �           �   s       ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f �M     �   r   t   �      4        H_0 => to_bitvector(unsigned(16#6a09e667#)),5��    r                     M                     5�_�   �   �           �   s       ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f �M     �   r   t   �      ,        H_0 => to_bitvector((16#6a09e667#)),5��    r                     M                     5�_�   �   �           �   s   (    ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f �O     �   r   t   �      +        H_0 => to_bitvector(16#6a09e667#)),5��    r   (                  Y                     5�_�   �   �           �   s       ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f �d     �   r   t   �      *        H_0 => to_bitvector(16#6a09e667#),5��    r                     M                     5�_�   �   �           �   t       ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f �|     �   s   u   �              H_1 => 16#bb67ae85#,5��    s                     o                     5�_�   �   �           �   t   ,    ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f      �   s   u   �      -        H_1 => to_bitvector(32, 16#bb67ae85#,5��    s   ,                  �                     5�_�   �   �           �   u       ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f      �   t   v   �              H_2 => 16#3c6ef372#,5��    t                     �                     �    t   ,                  �                     5�_�   �   �           �   v       ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f      �   u   w   �              H_3 => 16#a54ff53a#,5��    u                     �                     �    u   ,                  �                     5�_�   �   �           �   w       ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f      �   v   x   �              H_4 => 16#510e527f#,5��    v                     �                     �    v   ,                                       5�_�   �   �           �   x       ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f      �   w   y   �              H_5 => 16#9b05688c#,5��    w                     +                     �    w   ,                  H                     5�_�   �   �           �   y       ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f      �   x   z   �              H_6 => 16#1f83d9ab#,5��    x                     Z                     �    x   ,                  w                     5�_�   �   �           �   z       ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f      �   y   {   �              H_7 => 16#5be0cd19#5��    y                     �                     5�_�   �   �           �   z   ,    ����                                                                                                                                                                                                                                                                                                                $                        !       v   !    f      �   y   {   �      ,        H_7 => to_bitvector(32, 16#5be0cd19#5��    y   ,                  �                     5�_�   �   �           �   e        ����                                                                                                                                                                                                                                                                                                                $           r          {          V   ,    f ®     �   e   g   �    5��    e                      �                     �    e                      �                     5�_�   �   �           �   f        ����                                                                                                                                                                                                                                                                                                                $           s          |          V   ,    f °     �   f   q   �    �   f   g   �    5��    f               
       �              �      5�_�   �   �           �   g       ����                                                                                                                                                                                                                                                                                                                $           }          �          V   ,    f ²     �   f   h   �          constant H : h_vector := (5��    f                    �                    5�_�   �   �           �   g       ����                                                                                                                                                                                                                                                                                                                $           }          �          V   ,    f ´     �   f   h   �          constant K : h_vector := (5��    f                    �                    5�_�   �   �           �   h        ����                                                                                                                                                                                                                                                                                                                $           h          n          V       f º     �   g   h          .        H_0 => to_bitvector(32, 16#6a09e667#),   .        H_1 => to_bitvector(32, 16#bb67ae85#),   .        H_2 => to_bitvector(32, 16#3c6ef372#),   .        H_3 => to_bitvector(32, 16#a54ff53a#),   .        H_4 => to_bitvector(32, 16#510e527f#),   .        H_5 => to_bitvector(32, 16#9b05688c#),   .        H_6 => to_bitvector(32, 16#1f83d9ab#),5��    g                      �      I              5�_�   �   �           �   h       ����                                                                                                                                                                                                                                                                                                                $           d          %          V       f ��     �   g   �   �    �   h   i   �    5��    g               @       �              �	      5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                $           h          �          V       f ��     �   �   �          -        H_7 => to_bitvector(32, 16#5be0cd19#)5��    �                      �      .               5�_�   �   �           �   h       ����                                                                                                                                                                                                                                                                                                                $           h          �          V       f ��     �   g   i   �    �   h   i   �    5��    g                      �              .       5�_�   �   �           �   i        ����                                                                                                                                                                                                                                                                                                                $           i          �          V       f ��     �   �   �          '        K_63 : bit_vector(31 downto 0);�   �   �          '        K_62 : bit_vector(31 downto 0);�   �   �          '        K_61 : bit_vector(31 downto 0);�   �   �          '        K_60 : bit_vector(31 downto 0);�   �   �          '        K_59 : bit_vector(31 downto 0);�   �   �          '        K_58 : bit_vector(31 downto 0);�   �   �          '        K_57 : bit_vector(31 downto 0);�   �   �          '        K_56 : bit_vector(31 downto 0);�   �   �          '        K_55 : bit_vector(31 downto 0);�   �   �          '        K_54 : bit_vector(31 downto 0);�   �   �          '        K_53 : bit_vector(31 downto 0);�   �   �          '        K_52 : bit_vector(31 downto 0);�   �   �          '        K_51 : bit_vector(31 downto 0);�   �   �          '        K_50 : bit_vector(31 downto 0);�   �   �          '        K_49 : bit_vector(31 downto 0);�   �   �          '        K_48 : bit_vector(31 downto 0);�   �   �          '        K_47 : bit_vector(31 downto 0);�   �   �          '        K_46 : bit_vector(31 downto 0);�   �   �          '        K_45 : bit_vector(31 downto 0);�   �   �          '        K_44 : bit_vector(31 downto 0);�   �   �          '        K_43 : bit_vector(31 downto 0);�   �   �          '        K_42 : bit_vector(31 downto 0);�   �   �          '        K_41 : bit_vector(31 downto 0);�   �   �          '        K_40 : bit_vector(31 downto 0);�   �   �          '        K_39 : bit_vector(31 downto 0);�   �   �          '        K_38 : bit_vector(31 downto 0);�   �   �          '        K_37 : bit_vector(31 downto 0);�   �   �          '        K_36 : bit_vector(31 downto 0);�   �   �          '        K_35 : bit_vector(31 downto 0);�   �   �          '        K_34 : bit_vector(31 downto 0);�   �   �          '        K_33 : bit_vector(31 downto 0);�   �   �          '        K_32 : bit_vector(31 downto 0);�   �   �          '        K_31 : bit_vector(31 downto 0);�   �   �          '        K_30 : bit_vector(31 downto 0);�   �   �          '        K_29 : bit_vector(31 downto 0);�   �   �          '        K_28 : bit_vector(31 downto 0);�   �   �          '        K_27 : bit_vector(31 downto 0);�   �   �          '        K_26 : bit_vector(31 downto 0);�   �   �          '        K_25 : bit_vector(31 downto 0);�   �   �          '        K_24 : bit_vector(31 downto 0);�      �          '        K_23 : bit_vector(31 downto 0);�   ~   �          '        K_22 : bit_vector(31 downto 0);�   }             '        K_21 : bit_vector(31 downto 0);�   |   ~          '        K_20 : bit_vector(31 downto 0);�   {   }          '        K_19 : bit_vector(31 downto 0);�   z   |          '        K_18 : bit_vector(31 downto 0);�   y   {          '        K_17 : bit_vector(31 downto 0);�   x   z          '        K_16 : bit_vector(31 downto 0);�   w   y          '        K_15 : bit_vector(31 downto 0);�   v   x          '        K_14 : bit_vector(31 downto 0);�   u   w          '        K_13 : bit_vector(31 downto 0);�   t   v          '        K_12 : bit_vector(31 downto 0);�   s   u          '        K_11 : bit_vector(31 downto 0);�   r   t          '        K_10 : bit_vector(31 downto 0);�   q   s          &        K_9 : bit_vector(31 downto 0);�   p   r          &        K_8 : bit_vector(31 downto 0);�   o   q          &        K_7 : bit_vector(31 downto 0);�   n   p          &        K_6 : bit_vector(31 downto 0);�   m   o          &        K_5 : bit_vector(31 downto 0);�   l   n          &        K_4 : bit_vector(31 downto 0);�   k   m          &        K_3 : bit_vector(31 downto 0);�   j   l          &        K_2 : bit_vector(31 downto 0);�   i   k          &        K_1 : bit_vector(31 downto 0);�   h   j   �      &        K_0 : bit_vector(31 downto 0);5��    h                                        �    i                    %                    �    j                    H                    �    k                    k                    �    l                    �                    �    m                    �                    �    n                    �                    �    o                    �                    �    p                                        �    q                    =                    �    r                    a                    �    s                    �                    �    t                    �                    �    u                    �                    �    v                    �                    �    w                                        �    x                    9                    �    y                    ]                    �    z                    �                    �    {                    �                    �    |                    �                    �    }                    �                    �    ~                                        �                        5                    �    �                    Y                    �    �                    }                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                                        �    �                    1                    �    �                    U                    �    �                    y                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    	                    �    �                    -                    �    �                    Q                    �    �                    u                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                                        �    �                    )                    �    �                    M                    �    �                    q                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                                        �    �                    %                    �    �                    I                    �    �                    m                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    !                    �    �                    E                    �    �                    i                    �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   �   #    ����                                                                                                                                                                                                                                                                                                                $           i          �          V       f �      �   �   �   �      #        K_63 => to_bitvector(32, ),5��    �   "                  �                     5�_�   �   �           �   i        ����                                                                                                                                                                                                                                                                                                                $           i   !       �   !       V   !    f �\     �   �   �          "        K_63 => to_bitvector(32, )�   �   �          #        K_62 => to_bitvector(32, ),�   �   �          #        K_61 => to_bitvector(32, ),�   �   �          #        K_60 => to_bitvector(32, ),�   �   �          #        K_59 => to_bitvector(32, ),�   �   �          #        K_58 => to_bitvector(32, ),�   �   �          #        K_57 => to_bitvector(32, ),�   �   �          #        K_56 => to_bitvector(32, ),�   �   �          #        K_55 => to_bitvector(32, ),�   �   �          #        K_54 => to_bitvector(32, ),�   �   �          #        K_53 => to_bitvector(32, ),�   �   �          #        K_52 => to_bitvector(32, ),�   �   �          #        K_51 => to_bitvector(32, ),�   �   �          #        K_50 => to_bitvector(32, ),�   �   �          #        K_49 => to_bitvector(32, ),�   �   �          #        K_48 => to_bitvector(32, ),�   �   �          #        K_47 => to_bitvector(32, ),�   �   �          #        K_46 => to_bitvector(32, ),�   �   �          #        K_45 => to_bitvector(32, ),�   �   �          #        K_44 => to_bitvector(32, ),�   �   �          #        K_43 => to_bitvector(32, ),�   �   �          #        K_42 => to_bitvector(32, ),�   �   �          #        K_41 => to_bitvector(32, ),�   �   �          #        K_40 => to_bitvector(32, ),�   �   �          #        K_39 => to_bitvector(32, ),�   �   �          #        K_38 => to_bitvector(32, ),�   �   �          #        K_37 => to_bitvector(32, ),�   �   �          #        K_36 => to_bitvector(32, ),�   �   �          #        K_35 => to_bitvector(32, ),�   �   �          #        K_34 => to_bitvector(32, ),�   �   �          #        K_33 => to_bitvector(32, ),�   �   �          #        K_32 => to_bitvector(32, ),�   �   �          #        K_31 => to_bitvector(32, ),�   �   �          #        K_30 => to_bitvector(32, ),�   �   �          #        K_29 => to_bitvector(32, ),�   �   �          #        K_28 => to_bitvector(32, ),�   �   �          #        K_27 => to_bitvector(32, ),�   �   �          #        K_26 => to_bitvector(32, ),�   �   �          #        K_25 => to_bitvector(32, ),�   �   �          #        K_24 => to_bitvector(32, ),�      �          #        K_23 => to_bitvector(32, ),�   ~   �          #        K_22 => to_bitvector(32, ),�   }             #        K_21 => to_bitvector(32, ),�   |   ~          #        K_20 => to_bitvector(32, ),�   {   }          #        K_19 => to_bitvector(32, ),�   z   |          #        K_18 => to_bitvector(32, ),�   y   {          #        K_17 => to_bitvector(32, ),�   x   z          #        K_16 => to_bitvector(32, ),�   w   y          #        K_15 => to_bitvector(32, ),�   v   x          #        K_14 => to_bitvector(32, ),�   u   w          #        K_13 => to_bitvector(32, ),�   t   v          #        K_12 => to_bitvector(32, ),�   s   u          #        K_11 => to_bitvector(32, ),�   r   t          #        K_10 => to_bitvector(32, ),�   q   s          "        K_9 => to_bitvector(32, ),�   p   r          "        K_8 => to_bitvector(32, ),�   o   q          "        K_7 => to_bitvector(32, ),�   n   p          "        K_6 => to_bitvector(32, ),�   m   o          "        K_5 => to_bitvector(32, ),�   l   n          "        K_4 => to_bitvector(32, ),�   k   m          "        K_3 => to_bitvector(32, ),�   j   l          "        K_2 => to_bitvector(32, ),�   i   k          "        K_1 => to_bitvector(32, ),�   h   j   �      "        K_0 => to_bitvector(32, ),5��    h                                        �    i                    :                    �    j                    a                    �    k                    �                    �    l                    �                    �    m                    �                    �    n                    �                    �    o                    $                    �    p                    K                    �    q                    r                    �    r                    �                    �    s                    �                    �    t                    �                    �    u                                        �    v                    :                    �    w                    b                    �    x                    �                    �    y                    �                    �    z                    �                    �    {                                        �    |                    *                    �    }                    R                    �    ~                    z                    �                        �                    �    �                    �                    �    �                    �                    �    �                                        �    �                    B                    �    �                    j                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    
                    �    �                    2                    �    �                    Z                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    "                    �    �                    J                    �    �                    r                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                                        �    �                    :                    �    �                    b                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                                        �    �                    *                    �    �                    R                    �    �                    z                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                                        �    �                    B                    �    �                    j                    �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   h       ����                                                                                                                                                                                                                                                                                                                $           i   !       �   !       V   !    f �d     �   g   h          -        H_7 => to_bitvector(32, 16#5be0cd19#)5��    g                      �      .               5�_�   �   �           �   h       ����                                                                                                                                                                                                                                                                                                                $           h   !       �   !       V   !    f �x     �   g   p   �          �   h   i   �    �   g   i   �    5��    g                      �              	       �    g                     �                    �    g                 G   �              ?      5�_�   �   �           �   h       ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f �{     �   g   i   �      K    428a2f98 71374491 b5c0fbcf e9b5dba5 3956c25b 59f111f1 923f82a4 ab1c5ed55��    g                      �                     5�_�   �   �           �   h        ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f É     �   g   i   �      G428a2f98 71374491 b5c0fbcf e9b5dba5 3956c25b 59f111f1 923f82a4 ab1c5ed55��    g           G           �      G               5�_�   �   �           �   p   "    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f Ñ     �   o   q   �      &        K_0 => to_bitvector(32, 16##),�   p   q   �    5��    o   #               G   �              G       5�_�   �   �           �   p   +    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f â     �   o   q   �      m        K_0 => to_bitvector(32, 16#428a2f98 71374491 b5c0fbcf e9b5dba5 3956c25b 59f111f1 923f82a4 ab1c5ed5#),5��    o   +                  �                     5�_�   �   �           �   p   +    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f å     �   o   q   �      l        K_0 => to_bitvector(32, 16#428a2f9871374491 b5c0fbcf e9b5dba5 3956c25b 59f111f1 923f82a4 ab1c5ed5#),5��    o   +       >           �      >               5�_�   �   �           �   q   "    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ì     �   p   r   �      &        K_1 => to_bitvector(32, 16##),�   q   r   �    5��    p   #               >                 >       5�_�   �   �           �   q   +    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ó     �   q   s   �      &        K_2 => to_bitvector(32, 16##),�   r   s   �    �   p   r   �      d        K_1 => to_bitvector(32, 16#71374491 b5c0fbcf e9b5dba5 3956c25b 59f111f1 923f82a4 ab1c5ed5#),5��    p   +                                       �    p   +       5                 5               �    q   #               5   B              5       5�_�   �   �           �   r   +    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ÿ     �   v   x   �      &        K_7 => to_bitvector(32, 16##),�   w   x   �    �   u   w   �      &        K_6 => to_bitvector(32, 16##),�   v   w   �    �   t   v   �      &        K_5 => to_bitvector(32, 16##),�   u   v   �    �   s   u   �      &        K_4 => to_bitvector(32, 16##),�   t   u   �    �   r   t   �      &        K_3 => to_bitvector(32, 16##),�   s   t   �    �   q   s   �      [        K_2 => to_bitvector(32, 16#b5c0fbcf e9b5dba5 3956c25b 59f111f1 923f82a4 ab1c5ed5#),5��    q   +                  J                     �    q   +       ,           J      ,               �    r   #               ,   q              ,       �    r   +       $           y      $               �    s   #               #   �              #       �    s   +                  �                     �    t   #                  �                     �    t   +                  �                     �    u   #                  �                     �    u   +       	                 	               �    v   #                  -                     5�_�   �   �           �   i        ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ��     �   h   j   �      Gd807aa98 12835b01 243185be 550c7dc3 72be5d74 80deb1fe 9bdc06a7 c19bf1745��    h           G           �      G               5�_�   �   �           �   x   "    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ��     �   w   y   �      &        K_8 => to_bitvector(32, 16##),�   x   y   �    5��    w   #               G                 G       5�_�   �   �           �   x   +    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ��     �   ~   �   �      '        K_15 => to_bitvector(32, 16##),�      �   �    �   }      �      '        K_14 => to_bitvector(32, 16##),�   ~      �    �   |   ~   �      '        K_13 => to_bitvector(32, 16##),�   }   ~   �    �   {   }   �      '        K_12 => to_bitvector(32, 16##),�   |   }   �    �   z   |   �      '        K_11 => to_bitvector(32, 16##),�   {   |   �    �   y   {   �      '        K_10 => to_bitvector(32, 16##),�   z   {   �    �   x   z   �      &        K_9 => to_bitvector(32, 16##),�   y   z   �    �   w   y   �      m        K_8 => to_bitvector(32, 16#d807aa98 12835b01 243185be 550c7dc3 72be5d74 80deb1fe 9bdc06a7 c19bf174#),5��    w   +                                       �    w   +       >                 >               �    x   #               >   D              >       �    x   +       6           L      6               �    y   $               5   t              5       �    y   ,       -           |      -               �    z   $               ,   �              ,       �    z   ,       $           �      $               �    {   $               #   �              #       �    {   ,                  �                     �    |   $                                       �    |   ,                                       �    }   $                  4                     �    }   ,       	           <      	               �    ~   $                  d                     5�_�   �   �           �   j        ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ��     �   i   k   �      Ge49b69c1 efbe4786 0fc19dc6 240ca1cc 2de92c6f 4a7484aa 5cb0a9dc 76f988da5��    i           G           �      G               5�_�   �   �           �   �   #    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ��     �      �   �      '        K_16 => to_bitvector(32, 16##),�   �   �   �    5��       $               G   M              G       5�_�   �   �           �   �   ,    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ��     �   �   �   �      '        K_23 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_22 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_21 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_20 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_19 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_18 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_17 => to_bitvector(32, 16##),�   �   �   �    �      �   �      n        K_16 => to_bitvector(32, 16#e49b69c1 efbe4786 0fc19dc6 240ca1cc 2de92c6f 4a7484aa 5cb0a9dc 76f988da#),5��       ,                  U                     �       ,       >           U      >               �    �   $               >   }              >       �    �   ,       6           �      6               �    �   $               5   �              5       �    �   ,       -           �      -               �    �   $               ,   �              ,       �    �   ,       $           �      $               �    �   $               #                 #       �    �   ,                                       �    �   $                  =                     �    �   ,                  E                     �    �   $                  m                     �    �   ,       	           u      	               �    �   $                  �                     5�_�   �   �           �   k        ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ��     �   j   l   �      G983e5152 a831c66d b00327c8 bf597fc7 c6e00bf3 d5a79147 06ca6351 142929675��    j           G           �      G               5�_�   �   �           �   �   #    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ��     �   �   �   �      '        K_24 => to_bitvector(32, 16##),�   �   �   �    5��    �   $               G   �              G       5�_�   �   �           �   �   ,    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ��     �   �   �   �      '        K_31 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_30 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_29 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_28 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_27 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_26 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_25 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      n        K_24 => to_bitvector(32, 16#983e5152 a831c66d b00327c8 bf597fc7 c6e00bf3 d5a79147 06ca6351 14292967#),5��    �   ,                  �                     �    �   ,       >           �      >               �    �   $               >   �              >       �    �   ,       6           �      6               �    �   $               5   �              5       �    �   ,       -           �      -               �    �   $               ,                 ,       �    �   ,       $                 $               �    �   $               #   F              #       �    �   ,                  N                     �    �   $                  v                     �    �   ,                  ~                     �    �   $                  �                     �    �   ,       	           �      	               �    �   $                  �                     5�_�   �   �           �   l        ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ��     �   k   m   �      G27b70a85 2e1b2138 4d2c6dfc 53380d13 650a7354 766a0abb 81c2c92e 92722c855��    k           G           �      G               5�_�   �   �           �   �   #    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ��     �   �   �   �      '        K_32 => to_bitvector(32, 16##),�   �   �   �    5��    �   $               G   �              G       5�_�   �   �           �   �   ,    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ��     �   �   �   �      '        K_39 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_38 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_37 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_36 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_35 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_34 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_33 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      n        K_32 => to_bitvector(32, 16#27b70a85 2e1b2138 4d2c6dfc 53380d13 650a7354 766a0abb 81c2c92e 92722c85#),5��    �   ,                  �                     �    �   ,       >           �      >               �    �   $               >   �              >       �    �   ,       6           �      6               �    �   $               5                 5       �    �   ,       -           '      -               �    �   $               ,   O              ,       �    �   ,       $           W      $               �    �   $               #                 #       �    �   ,                  �                     �    �   $                  �                     �    �   ,                  �                     �    �   $                  �                     �    �   ,       	           �      	               �    �   $                                       5�_�   �   �           �   m        ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f ��     �   l   n   �      Ga2bfe8a1 a81a664b c24b8b70 c76c51a3 d192e819 d6990624 f40e3585 106aa0705��    l           G           �      G               5�_�   �   �           �   �   #    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f �     �   �   �   �      '        K_40 => to_bitvector(32, 16##),�   �   �   �    5��    �   $               G   �              G       5�_�   �   �           �   �   ,    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f �     �   �   �   �      '        K_47 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_46 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_45 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_44 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_43 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_42 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_41 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      n        K_40 => to_bitvector(32, 16#a2bfe8a1 a81a664b c24b8b70 c76c51a3 d192e819 d6990624 f40e3585 106aa070#),5��    �   ,                                        �    �   ,       >                  >               �    �   $               >   (              >       �    �   ,       6           0      6               �    �   $               5   X              5       �    �   ,       -           `      -               �    �   $               ,   �              ,       �    �   ,       $           �      $               �    �   $               #   �              #       �    �   ,                  �                     �    �   $                  �                     �    �   ,                  �                     �    �   $                                       �    �   ,       	                  	               �    �   $                  H                     5�_�   �   �   �       �   n        ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f �     �   m   o   �      G19a4c116 1e376c08 2748774c 34b0bcb5 391c0cb3 4ed8aa4a 5b9cca4f 682e6ff35��    m           G           �      G               5�_�   �   �           �   �   #    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f �     �   �   �   �      '        K_48 => to_bitvector(32, 16##),�   �   �   �    5��    �   $               G   1              G       5�_�   �   �           �   �   ,    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f �     �   �   �   �      '        K_55 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_54 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_53 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_52 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_51 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_50 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_49 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      n        K_48 => to_bitvector(32, 16#19a4c116 1e376c08 2748774c 34b0bcb5 391c0cb3 4ed8aa4a 5b9cca4f 682e6ff3#),5��    �   ,                  9                     �    �   ,       >           9      >               �    �   $               >   a              >       �    �   ,       6           i      6               �    �   $               5   �              5       �    �   ,       -           �      -               �    �   $               ,   �              ,       �    �   ,       $           �      $               �    �   $               #   �              #       �    �   ,                  �                     �    �   $                  !                     �    �   ,                  )                     �    �   $                  Q                     �    �   ,       	           Y      	               �    �   $                  �                     5�_�   �   �           �   o        ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f �     �   n   p   �      G748f82ee 78a5636f 84c87814 8cc70208 90befffa a4506ceb bef9a3f7 c67178f25��    n           G           �      G               5�_�   �   �           �   �   #    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f �#     �   �   �   �      '        K_56 => to_bitvector(32, 16##),�   �   �   �    5��    �   $               G   j              G       5�_�   �   �           �   �   ,    ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f �*     �   �   �   �      &        K_63 => to_bitvector(32, 16##)�   �   �   �    �   �   �   �      '        K_62 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_61 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_60 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_59 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_58 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      '        K_57 => to_bitvector(32, 16##),�   �   �   �    �   �   �   �      n        K_56 => to_bitvector(32, 16#748f82ee 78a5636f 84c87814 8cc70208 90befffa a4506ceb bef9a3f7 c67178f2#),5��    �   ,                  r                     �    �   ,       >           r      >               �    �   $               >   �              >       �    �   ,       6           �      6               �    �   $               5   �              5       �    �   ,       -           �      -               �    �   $               ,   �              ,       �    �   ,       $                 $               �    �   $               #   *              #       �    �   ,                  2                     �    �   $                  Z                     �    �   ,                  b                     �    �   $                  �                     �    �   ,       	           �      	               �    �   $                  �                     5�_�   �   �           �   h        ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f �.     �   g   h                                       5��    g                      �                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                $           h   !       �   !       V   !    f �i     �          �    5��                                                  5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                %           i   !       �   !       V   !    f �j     �          �       �         �    �          �    5��                                                  �                    
                      K      5�_�   �   �           �      	    ����                                                                                                                                                                                                                                                                                                                0           t   !       �   !       V   !    f �o     �         �      use IEEE.NUMERIC_STD.ALL;5��       	                 4                     �       
                  5                      �       	                 4                     �       	                 4                     �       	                 4                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                0           t   !       �   !       V   !    f �x     �      	   �      ?        reset : in bit;                          -- Reset input5��                        �                     5�_�   �   �           �   	       ����                                                                                                                                                                                                                                                                                                                0           t   !       �   !       V   !    f ń     �      
   �      F        count : out bit_vector(2 downto 0)       -- 3-bit count output5��                                            5�_�   �   �           �   	       ����                                                                                                                                                                                                                                                                                                                0           t   !       �   !       V   !    f ŋ     �      
   �      F        count : out bit_vector(7 downto 0)       -- 3-bit count output5��                                            5�_�   �   �           �   	   4    ����                                                                                                                                                                                                                                                                                                                0           t   !       �   !       V   !    f ŏ     �      
   �      F        count : out bit_vector(5 downto 0)       -- 3-bit count output5��       4                                     5�_�   �   �           �   	   F    ����                                                                                                                                                                                                                                                                                                                0           t   !       �   !       V   !    f ő     �      
   �      F        count : out bit_vector(5 downto 0)       -- 6-bit count output5��       F                  .                     5�_�   �   �           �   	   G    ����                                                                                                                                                                                                                                                                                                                0           t   !       �   !       V   !    f Œ     �      
   �      G        count : out bit_vector(5 downto 0)       -- 6-bit count output 5��       G                  /                     5�_�   �   �           �   	   H    ����                                                                                                                                                                                                                                                                                                                0           t   !       �   !       V   !    f œ     �      
   �      I        count : out bit_vector(5 downto 0)       -- 6-bit count output ()5��       H                  0                     �       I                 1                    5�_�   �   �           �   	   J    ����                                                                                                                                                                                                                                                                                                                0           t   !       �   !       V   !    f ŕ     �      
   �      K        count : out bit_vector(5 downto 0)       -- 6-bit count output (64)5��       J                  2                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                0           t   !       �   !       V   !    f ŝ     �         �      entity Binary_Counter is5��                        M                     �                        Q                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                0           t   !       �   !       V   !    f Ť     �         �      entity couter is5��                         S                      5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                0           t   !       �   !       V   !    f Ũ     �   
      �      end Binary_Counter;5��    
                    B                    �    
                     F                     �    
                    E                    �    
                    E                    �    
                     E                     �    
                     D                     �    
                     C                     �    
                    B                    �    
                    B                    �    
                    B                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                0           t   !       �   !       V   !    f Ű     �         �      end architecture �         �      architecture rtl of  is�         �          �         �      arch�         �       �         �    5��                          O                     �                          O                     �                          P                     �                         S                     �                         R                     �                         Q                     �                         P                    �                         P                    �                         P                    �                         P                    �                        d                     �                          |                      �                        |                     �                         �                     �                      
   d              
       �                         �                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                8                               v       f Ŷ     �         �      !architecture rtl of multisteps is5��              
          d      
              5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                8                               v       f ��     �   
      �      end couter_6bit;5��    
                     E                     5�_�   �   �           �      
    ����                                                                                                                                                                                                                                                                                                                8                               v       f ��     �         �      entity couter_6bit is5��       
                  P                      5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                8                               v       f ��     �         �          5��                         z                     �                         {                     �                        z                    �                         {                     �                        z                    �                        z                    �                        z                    �                        z                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                8                               v       f ��     �         �          signed(7 downto 0)5��                        z                    �                        {                    �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    �                        �                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                8                               v       f ��     �         �      (    signal counter: unsigned(7 downto 0)5��                        �                    5�_�   �   �           �      (    ����                                                                                                                                                                                                                                                                                                                8                               v       f ��     �         �      (    signal counter: unsigned(5 downto 0)5��       (                  �                     �       )                 �                     �                         �                     �                         �                     �                         �                     �                          �                     5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                9                               v       f ��     �         �          end process �         �              �         �          5��                         �                     �                         �                     �                         �                     �                        �                    �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �       
                  �                     �       	                  �                     �                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �       
                  �                     �       	                  �                     �                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �       
                  �                     �       	                  �                     �                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �       
                  �                     �       	                  �                     �                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    �                     #   �             #       �       '                 �                     �                          �                      �                        �                     �                      
   �              
       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                <                               v       f �7     �         �    �         �          end process proc_name;�         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �      (    proc_name: process(sensitivity_list)5��              	          �      	              �              	          �      	              �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �       	                  �                     �                        �                    �       
                  �                     �                        �                    �                         �                     �                        �                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                <              %                 v       f �C     �         �              �         �      '    counting: process(sensitivity_list)5��                        �                    �                         �                     �                        �                    �                        �                    �                        �                    �                         �                     �                        �                    �                        �                    �                        �                    �                         �                     �                        �                    �                         �                     �                        �                    �                        �                    �                        �                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                <              %                 v       f �Z     �         �              if rst = 5��                         �                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                <              %                 v       f �[     �         �              if rst = ''5��                         �                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                <              %                 v       f �]     �         �                  counter�         �              if rst = '1'5��                         �                     �                         �                     �                        �              	       �                         �                    �                         �                     �                         �                     �                         �                     �                        �                    �                                              �                                              �                                              �                                              �                                              �                                              �                                              �                                               �                         �                     �                         �                     �                         �                     �                        �                    �                                              �                                              �                                              �                                               �                         �                     �                         �                     �                         �                     �                        �                    �                                              �                                              �                                               �                         �                     �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    �                         	                     �                                              �                                            �                         	                     �                                              �                                            �                                            �                                            �                                            5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                =              %                 v       f �r     �         �      $            counter => others => '0'5��                                              5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                =              %                 v       f �s     �         �      #            counter = others => '0'5��                                              5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                =              %                 v       f �u     �         �      $            counter <= others => '0'5��                                              5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                =              %                 v       f �~     �         �      %            counter <= (others => '0'5��                         �      &       '       5�_�   �   �           �      $    ����                                                                                                                                                                                                                                                                                                                =              %                 v       f Ɓ     �         �      &            counter <= (others => '0)'5��       $                                       5�_�   �   �           �      $    ����                                                                                                                                                                                                                                                                                                                =              %                 v       f Ɓ     �         �      %            counter <= (others => '0'�         �    5��       %                                       5�_�   �   �           �      &    ����                                                                                                                                                                                                                                                                                                                =              %                 v       f Ƃ     �         �      &            counter <= (others => '0')5��       &                                       5�_�   �   �           �      &    ����                                                                                                                                                                                                                                                                                                                =              %                 v       f Ƅ     �         �                  �         �    5��                                               �                         $                     �                        &                    �                                             �                         $                     �                         %                     �                         $                     �                         #                     �       
                  "                     �       	                 !                    �       
                 "                    �                         #                     �       
                 "                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                >              %                 v       f Ƙ     �         �              elsif rising_edge5��                         1                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                >              %                 v       f ƛ     �         �              elsif rising_edge()5��                         2                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                >              %                 v       f Ɯ     �         �                  counter�         �              elsif rising_edge(clk)5��                         6                     �                        7                    �                        7                    �                        7                    �       #                 ;              	       �                         <                    �                         K                     �                         J                     �                         I                     �                        H                    �                        H                    �                     
   H             
       �                        Q                    �                        U                    �                         W                     �                         V                     �                         U                     �                         T                     �                        S                    �                         W                     �                         V                     �                         U                     �                         T                     �                        S                    �                         Y                     �                         X                     �                         W                     �                         V                     �                         U                     �                         T                     �                        S                    �                        S                    �                        S                    �       #                 _                     �                         l                     �                         `                    �                         l                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                @              %                 v       f ƾ     �         �          count <= bit_vector�         �          �         �    5��                          �                     �                          �                     �                         �                     �                         �                     �                         �                     �                        �                    �                        �                    �                         �                     �                        �                    �                         �                     �                         �                     �                         �                     �                     
   �             
       �              
          �      
              �                     
   �             
       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                B              %                 v       f ��     �         �          count <= bit_vector5��                         �                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                B              %                 v       f ��     �         �          count <= bit_vector()5��                         �                     �                        �                    �                        �                    �                        �                    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                B              %                 v       f ��    �         �           count <= bit_vector(counter)5��                          �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                B           .   	       7   	       V   	    f�=     �   �   �   �      .        K_0 => to_bitvector(32, 16#428a2f98#),5��    �          	          �      	              5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                B           .   	       7   	       V   	    f�M     �   �   �   �      +        K_0 => to_signed(32, 16#428a2f98#),5��    �                     �                     �    �                     �                     5�_�   �   �           �   �   +    ����                                                                                                                                                                                                                                                                                                                B           .   	       7   	       V   	    f�R     �   �   �   �      ,        K_0 => (to_signed(32, 16#428a2f98#),5��    �   +                  �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                B           .   	       7   	       V   	    f�Z     �   �   �   �      -        K_0 => (to_signed(32, 16#428a2f98#)),5��    �                     �                     �    �                     �                     �    �                    �                    �    �                     �                     �    �                 
   �             
       �    �          
       
   �      
       
       �    �          
          �      
              �    �                 
   �             
       5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                B           �          �          V       f̋     �   �   �          .        K_63 => to_bitvector(32, 16#c67178f2#)�   �   �          /        K_62 => to_bitvector(32, 16#bef9a3f7#),�   �   �          /        K_61 => to_bitvector(32, 16#a4506ceb#),�   �   �          /        K_60 => to_bitvector(32, 16#90befffa#),�   �   �          /        K_59 => to_bitvector(32, 16#8cc70208#),�   �   �          /        K_58 => to_bitvector(32, 16#84c87814#),�   �   �          /        K_57 => to_bitvector(32, 16#78a5636f#),�   �   �          /        K_56 => to_bitvector(32, 16#748f82ee#),�   �   �          /        K_55 => to_bitvector(32, 16#682e6ff3#),�   �   �          /        K_54 => to_bitvector(32, 16#5b9cca4f#),�   �   �          /        K_53 => to_bitvector(32, 16#4ed8aa4a#),�   �   �          /        K_52 => to_bitvector(32, 16#391c0cb3#),�   �   �          /        K_51 => to_bitvector(32, 16#34b0bcb5#),�   �   �          /        K_50 => to_bitvector(32, 16#2748774c#),�   �   �          /        K_49 => to_bitvector(32, 16#1e376c08#),�   �   �          /        K_48 => to_bitvector(32, 16#19a4c116#),�   �   �          /        K_47 => to_bitvector(32, 16#106aa070#),�   �   �          /        K_46 => to_bitvector(32, 16#f40e3585#),�   �   �          /        K_45 => to_bitvector(32, 16#d6990624#),�   �   �          /        K_44 => to_bitvector(32, 16#d192e819#),�   �   �          /        K_43 => to_bitvector(32, 16#c76c51a3#),�   �   �          /        K_42 => to_bitvector(32, 16#c24b8b70#),�   �   �          /        K_41 => to_bitvector(32, 16#a81a664b#),�   �   �          /        K_40 => to_bitvector(32, 16#a2bfe8a1#),�   �   �          /        K_39 => to_bitvector(32, 16#92722c85#),�   �   �          /        K_38 => to_bitvector(32, 16#81c2c92e#),�   �   �          /        K_37 => to_bitvector(32, 16#766a0abb#),�   �   �          /        K_36 => to_bitvector(32, 16#650a7354#),�   �   �          /        K_35 => to_bitvector(32, 16#53380d13#),�   �   �          /        K_34 => to_bitvector(32, 16#4d2c6dfc#),�   �   �          /        K_33 => to_bitvector(32, 16#2e1b2138#),�   �   �          /        K_32 => to_bitvector(32, 16#27b70a85#),�   �   �          /        K_31 => to_bitvector(32, 16#14292967#),�   �   �          /        K_30 => to_bitvector(32, 16#06ca6351#),�   �   �          /        K_29 => to_bitvector(32, 16#d5a79147#),�   �   �          /        K_28 => to_bitvector(32, 16#c6e00bf3#),�   �   �          /        K_27 => to_bitvector(32, 16#bf597fc7#),�   �   �          /        K_26 => to_bitvector(32, 16#b00327c8#),�   �   �          /        K_25 => to_bitvector(32, 16#a831c66d#),�   �   �          /        K_24 => to_bitvector(32, 16#983e5152#),�   �   �          /        K_23 => to_bitvector(32, 16#76f988da#),�   �   �          /        K_22 => to_bitvector(32, 16#5cb0a9dc#),�   �   �          /        K_21 => to_bitvector(32, 16#4a7484aa#),�   �   �          /        K_20 => to_bitvector(32, 16#2de92c6f#),�   �   �          /        K_19 => to_bitvector(32, 16#240ca1cc#),�   �   �          /        K_18 => to_bitvector(32, 16#0fc19dc6#),�   �   �          /        K_17 => to_bitvector(32, 16#efbe4786#),�   �   �          /        K_16 => to_bitvector(32, 16#e49b69c1#),�   �   �          /        K_15 => to_bitvector(32, 16#c19bf174#),�   �   �          /        K_14 => to_bitvector(32, 16#9bdc06a7#),�   �   �          /        K_13 => to_bitvector(32, 16#80deb1fe#),�   �   �          /        K_12 => to_bitvector(32, 16#72be5d74#),�   �   �          /        K_11 => to_bitvector(32, 16#550c7dc3#),�   �   �          /        K_10 => to_bitvector(32, 16#243185be#),�   �   �          .        K_9 => to_bitvector(32, 16#12835b01#),�   �   �          .        K_8 => to_bitvector(32, 16#d807aa98#),�   �   �          .        K_7 => to_bitvector(32, 16#ab1c5ed5#),�   �   �          .        K_6 => to_bitvector(32, 16#923f82a4#),�   �   �          .        K_5 => to_bitvector(32, 16#59f111f1#),�   �   �          .        K_4 => to_bitvector(32, 16#3956c25b#),�   �   �          .        K_3 => to_bitvector(32, 16#e9b5dba5#),�   �   �          .        K_2 => to_bitvector(32, 16#b5c0fbcf#),�   �   �   �      .        K_1 => to_bitvector(32, 16#71374491#),5��    �                    �                    �    �                                        �    �                    F                    �    �                    }                    �    �                    �                    �    �                    �                    �    �                    "                    �    �                    Y                    �    �                    �                    �    �                    �                    �    �                                         �    �                    8                    �    �                    p                    �    �                    �                    �    �                    �                    �    �                                        �    �                    P                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    0                    �    �                    h                    �    �                    �                    �    �                    �                    �    �                                        �    �                    H                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    (                    �    �                    `                    �    �                    �                    �    �                    �                    �    �                                        �    �                    @                    �    �                    x                    �    �                    �                    �    �                    �                    �    �                                         �    �                    X                    �    �                    �                    �    �                    �                    �    �                                         �    �                    8                    �    �                    p                    �    �                    �                    �    �                    �                    �    �                                        �    �                    P                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    0                    �    �                    h                    �    �                    �                    �    �                    �                    �    �                                        �    �                    H                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    (                    �    �                    `                    5�_�   �   �           �   �   5    ����                                                                                                                                                                                                                                                                                                                B           �   5       �   5          5    f̕    �   �   �   �   >   6        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#),   6        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#),   6        K_4 => bit_vector(to_signed(32, 16#3956c25b#),   6        K_5 => bit_vector(to_signed(32, 16#59f111f1#),   6        K_6 => bit_vector(to_signed(32, 16#923f82a4#),   6        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#),   6        K_8 => bit_vector(to_signed(32, 16#d807aa98#),   6        K_9 => bit_vector(to_signed(32, 16#12835b01#),   7        K_10 => bit_vector(to_signed(32, 16#243185be#),   7        K_11 => bit_vector(to_signed(32, 16#550c7dc3#),   7        K_12 => bit_vector(to_signed(32, 16#72be5d74#),   7        K_13 => bit_vector(to_signed(32, 16#80deb1fe#),   7        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#),   7        K_15 => bit_vector(to_signed(32, 16#c19bf174#),   7        K_16 => bit_vector(to_signed(32, 16#e49b69c1#),   7        K_17 => bit_vector(to_signed(32, 16#efbe4786#),   7        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#),   7        K_19 => bit_vector(to_signed(32, 16#240ca1cc#),   7        K_20 => bit_vector(to_signed(32, 16#2de92c6f#),   7        K_21 => bit_vector(to_signed(32, 16#4a7484aa#),   7        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#),   7        K_23 => bit_vector(to_signed(32, 16#76f988da#),   7        K_24 => bit_vector(to_signed(32, 16#983e5152#),   7        K_25 => bit_vector(to_signed(32, 16#a831c66d#),   7        K_26 => bit_vector(to_signed(32, 16#b00327c8#),   7        K_27 => bit_vector(to_signed(32, 16#bf597fc7#),   7        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#),   7        K_29 => bit_vector(to_signed(32, 16#d5a79147#),   7        K_30 => bit_vector(to_signed(32, 16#06ca6351#),   7        K_31 => bit_vector(to_signed(32, 16#14292967#),   7        K_32 => bit_vector(to_signed(32, 16#27b70a85#),   7        K_33 => bit_vector(to_signed(32, 16#2e1b2138#),   7        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#),   7        K_35 => bit_vector(to_signed(32, 16#53380d13#),   7        K_36 => bit_vector(to_signed(32, 16#650a7354#),   7        K_37 => bit_vector(to_signed(32, 16#766a0abb#),   7        K_38 => bit_vector(to_signed(32, 16#81c2c92e#),   7        K_39 => bit_vector(to_signed(32, 16#92722c85#),   7        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#),   7        K_41 => bit_vector(to_signed(32, 16#a81a664b#),   7        K_42 => bit_vector(to_signed(32, 16#c24b8b70#),   7        K_43 => bit_vector(to_signed(32, 16#c76c51a3#),   7        K_44 => bit_vector(to_signed(32, 16#d192e819#),   7        K_45 => bit_vector(to_signed(32, 16#d6990624#),   7        K_46 => bit_vector(to_signed(32, 16#f40e3585#),   7        K_47 => bit_vector(to_signed(32, 16#106aa070#),   7        K_48 => bit_vector(to_signed(32, 16#19a4c116#),   7        K_49 => bit_vector(to_signed(32, 16#1e376c08#),   7        K_50 => bit_vector(to_signed(32, 16#2748774c#),   7        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#),   7        K_52 => bit_vector(to_signed(32, 16#391c0cb3#),   7        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#),   7        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#),   7        K_55 => bit_vector(to_signed(32, 16#682e6ff3#),   7        K_56 => bit_vector(to_signed(32, 16#748f82ee#),   7        K_57 => bit_vector(to_signed(32, 16#78a5636f#),   7        K_58 => bit_vector(to_signed(32, 16#84c87814#),   7        K_59 => bit_vector(to_signed(32, 16#8cc70208#),   7        K_60 => bit_vector(to_signed(32, 16#90befffa#),   7        K_61 => bit_vector(to_signed(32, 16#a4506ceb#),   7        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#),   6        K_63 => bit_vector(to_signed(32, 16#c67178f2#)�   �   �   �      6        K_1 => bit_vector(to_signed(32, 16#71374491#),5��    �   5                  �                     �    �   5                  6                     �    �   5                  n                     �    �   5                  �                     �    �   5                  �                     �    �   5                                       �    �   5                  N                     �    �   5                  �                     �    �   5                  �                     �    �   5                  �                     �    �   5                  /                     �    �   5                  h                     �    �   5                  �                     �    �   5                  �                     �    �   5                                       �    �   5                  L                     �    �   5                  �                     �    �   5                  �                     �    �   5                  �                     �    �   5                  0                     �    �   5                  i                     �    �   5                  �                     �    �   5                  �                     �    �   5                                       �    �   5                  M                     �    �   5                  �                     �    �   5                  �                     �    �   5                  �                     �    �   5                  1                     �    �   5                  j                     �    �   5                  �                     �    �   5                  �                     �    �   5                                       �    �   5                  N                     �    �   5                  �                     �    �   5                  �                     �    �   5                  �                     �    �   5                  2                     �    �   5                  k                     �    �   5                  �                     �    �   5                  �                     �    �   5                                       �    �   5                  O                     �    �   5                  �                     �    �   5                  �                     �    �   5                  �                     �    �   5                  3                     �    �   5                  l                     �    �   5                  �                     �    �   5                  �                     �    �   5                                       �    �   5                  P                     �    �   5                  �                     �    �   5                  �                     �    �   5                  �                     �    �   5                  4                     �    �   5                  m                     �    �   5                  �                     �    �   5                  �                     �    �   5                                       �    �   5                  Q                     �    �   5                  �                     �    �   5                  �                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                B           �   )       �   )       V   )    f�(     �   �   �          -        H_7 => to_bitvector(32, 16#5be0cd19#)�   �   �          .        H_6 => to_bitvector(32, 16#1f83d9ab#),�   �   �          .        H_5 => to_bitvector(32, 16#9b05688c#),�   �   �          .        H_4 => to_bitvector(32, 16#510e527f#),�   �   �          .        H_3 => to_bitvector(32, 16#a54ff53a#),�   �   �          .        H_2 => to_bitvector(32, 16#3c6ef372#),�   �   �          .        H_1 => to_bitvector(32, 16#bb67ae85#),�   �   �   �      .        H_0 => to_bitvector(32, 16#6a09e667#),5��    �                    e                     �    �                    �                     �    �                    �                     �    �                    
!                    �    �                    A!                    �    �                    x!                    �    �                    �!                    �    �                    �!                    5�_�   �              �   �   5    ����                                                                                                                                                                                                                                                                                                                B           �   4       �   4          4    f�1    �   �   �   �      6        H_1 => bit_vector(to_signed(32, 16#bb67ae85#),   6        H_2 => bit_vector(to_signed(32, 16#3c6ef372#),   6        H_3 => bit_vector(to_signed(32, 16#a54ff53a#),   6        H_4 => bit_vector(to_signed(32, 16#510e527f#),   6        H_5 => bit_vector(to_signed(32, 16#9b05688c#),   6        H_6 => bit_vector(to_signed(32, 16#1f83d9ab#),   5        H_7 => bit_vector(to_signed(32, 16#5be0cd19#)�   �   �   �      6        H_0 => bit_vector(to_signed(32, 16#6a09e667#),5��    �   5                  �                      �    �   5                  �                      �    �   5                  �                      �    �   5                  3!                     �    �   5                  k!                     �    �   5                  �!                     �    �   5                  �!                     �    �   5                  "                     5�_�   �                .        ����                                                                                                                                                                                                                                                                                                                B           .   	       7   	       V   	    f�a     �   -   .       
   Kfunction to_bitvector(size : natural; value : integer) return bit_vector is   G    variable result : bit_vector(size - 1 downto 0) := (others => '0');   begin       for i in 0 to size - 1 loop   '        if (value and (2**i)) /= 0 then               result(i) := '1';           end if;       end loop;       return result;   end function;5��    -       
               �      ?              5�_�                  .        ����                                                                                                                                                                                                                                                                                                                8           .   	       .   	       V   	    f�a    �   -   .           5��    -                      �                     5�_�                      ����                                                                                                                                                                                                                                                                                                                7                               v       fv     �         �      #        elsif rising_edge(clk) then5��                         &                     5�_�                        ����                                                                                                                                                                                                                                                                                                                7                               v       fw     �         �              elsif  then5��                         &                     5�_�                        ����                                                                                                                                                                                                                                                                                                                7                               v       f|     �         �              elsif () then5��                         '                     �                        7                    5�_�                    #    ����                                                                                                                                                                                                                                                                                                                7                               v       f�     �         �      )        elsif (clk'event and clk = ) then5��       #                  ;                     5�_�                    $    ����                                                                                                                                                                                                                                                                                                                7                               v       f�   	 �         �      +        elsif (clk'event and clk = '') then5��       $                  <                     5�_�                 ,       ����                                                                                                                                                                                                                                                                                                                7                               V       f�     �   +   -   �      (architecture behavioral of multisteps is5��    +          
          �      
              5�_�                 �       ����                                                                                                                                                                                                                                                                                                                7                               V       f�     �   �   �   �      end architecture behavioral;5��    �          
          !      
              5�_�               5        ����                                                                                                                                                                                                                                                                                                                7                               V       f     �   5   >   �    �   5   6   �    5��    5                                           5�_�                 6       ����                                                                                                                                                                                                                                                                                                                ?                               V       f     �   5   7   �          component stepfun  is5��    5                                        �    5                                          �    5                                          �    5                                          �    5                                        �    5                                          �    5                                          �    5                                          �    5                                          �    5                                        �    5                                          �    5                                          �    5                                          �    5                                          �    5                                          �    5                                          �    5                                          �    5                                          �    5                                          �    5                                          �    5                                          �    5                                        �    5                                        �    5                                        5�_�                 8        ����                                                                                                                                                                                                                                                                                                                ?           8          :          V       f(   
 �   7   ;   �    �   8   9   �    �   7   8          D        	ai, bi, ci, di, ei, fi, gi, hi: in bit_vector(31 downto 0);   ,            kpw: in bit_vector(31 downto 0);   G            ao, bo, co, do, eo, fo, go, ho: out bit_vector(31 downto 0)5��    7                      .      �               �    7                      .              �       5�_�                 8       ����                                                                                                                                                                                                                                                                                                                ?           8          :                 fR    �   8   ;   �      =        rst : in bit;                          -- Reset input   Q        count : out bit_vector(5 downto 0)       -- 6-bit count output (64 steps)�   7   9   �      ?        clk : in bit;                            -- Clock input5��    7                     6                     �    8                     z                     �    9                     �                     5�_�                 �       ����                                                                                                                                                                                                                                                                                                                ?           8          :                 fn     �   �   �   �          �   �   �   �    5��    �                      "                     �    �                      "                     �    �                     "                     �    �                     "                     �    �                     "                     �    �                 
   "             
       5�_�                 �       ����                                                                                                                                                                                                                                                                                                                ?           8          :                 ft     �   �   �   �          �   �   �   �    5��    �                      "                     �    �                     "                     5�_�                 �       ����                                                                                                                                                                                                                                                                                                                ?           8          :                 f�     �   �   �   �          signal 5��    �                     ""                     �    �                    %"                    �    �                     &"                     �    �                    %"                    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                ?           8          :                 f�     �   �   �   �          signal clk: bit := 0;5��    �                     ."                     5�_�               �       ����                                                                                                                                                                                                                                                                                                                ?           8          :                 f�     �   �   �              signal clk: bit := ;5��    �                      "                     5�_�                 �        ����                                                                                                                                                                                                                                                                                                                ?           8          :                 f�     �   �   �   �          5��    �                     '"                     �    �                     ."                     �    �   
                  -"                     �    �   	                  ,"                     �    �                     +"                     �    �                     *"                     �    �                     )"                     �    �                     ("                     �    �                 
   '"             
       �    �                     0"                     �    �                     /"                     �    �                     ."                     �    �   
                  -"                     �    �   	                  ,"                     �    �                     +"                     �    �                     *"                     �    �                     )"                     �    �                     ("                     �    �                    '"                    �    �                     2"                     �    �                     1"                     �    �                     0"                     �    �                     /"                     �    �                     ."                     �    �   
                  -"                     �    �   	                  ,"                     �    �                     +"                     �    �                     *"                     �    �                     )"                     �    �                     ("                     �    �                    '"                    �    �                    '"                    �    �                    '"                    �    �                     2"                     �    �                     1"                     �    �                     0"                     �    �                     /"                     �    �                    ."                    5�_�                  �       ����                                                                                                                                                                                                                                                                                                                ?           8          :                 f�     �   �   �   �          counter: 5��    �                     0"                     �    �                     1"                     �    �                    0"                    �    �                    0"                    �    �                    0"                    �    �                     >"                     �    �                    ="                    �    �                    ="                    �    �                    ="                    5�_�    !              �   "    ����                                                                                                                                                                                                                                                                                                                ?           8          :                 f     �   �   �   �      "    counter: counter_6bit port map5��    �   "                  E"                     5�_�     "          !   �   #    ����                                                                                                                                                                                                                                                                                                                ?           8          :                 f     �   �   �   �      $    counter: counter_6bit port map()5��    �   "                  E"                     �    �   "                 E"                    5�_�  !  #          "   �   #    ����                                                                                                                                                                                                                                                                                                                ?           8          :                 f     �   �   �   �      #    counter: counter_6bit port map 5��    �   #                  F"                     5�_�  "  $          #   �   %    ����                                                                                                                                                                                                                                                                                                                ?           8          :                 f     �   �   �   �      %    counter: counter_6bit port map ()5��    �   %                  H"                     5�_�  #  %          $   �   $    ����                                                                                                                                                                                                                                                                                                                ?           8          :                 f$     �   �   �   �      &    counter: counter_6bit port map ();5��    �   $                  G"                     �    �   *                 M"                    5�_�  $  &          %   �       ����                                                                                                                                                                                                                                                                                                                ?           8          :                 f+     �   �   �   �          �   �   �   �    5��    �                      "                     �    �                     "                     �    �                    "                    �    �                     "                     �    �                     "                     �    �                     "                     �    �                    "                    �    �                    "                    �    �                    "                    �    �                     ."                     �    �                    -"                    �    �                     -"                     �    �                     ,"                     �    �                    +"                    �    �                     ."                     �    �                    -"                    �    �                    -"                    �    �                    -"                    �    �                    -"                    5�_�  %  '          &   �       ����                                                                                                                                                                                                                                                                                                                ?           �          �          v       fC     �   �   �   �      *    signal iteration: unsigned(7 downto 0)5��    �                    6"                    5�_�  &  (          '   �   *    ����                                                                                                                                                                                                                                                                                                                ?           �          �          v       fH     �   �   �   �      *    signal iteration: unsigned(5 downto 0)5��    �   *                  A"                     5�_�  '  )          (   �   .    ����                                                                                                                                                                                                                                                                                                                ?           �          �          v       fJ     �   �   �   �      .    signal iteration: unsigned(5 downto 0) := 5��    �   .                  E"                     5�_�  (  *          )   �   /    ����                                                                                                                                                                                                                                                                                                                ?           �          �          v       fK     �   �   �   �      0    signal iteration: unsigned(5 downto 0) := ""5��    �   /                  F"                     5�_�  )  +          *   �   6    ����                                                                                                                                                                                                                                                                                                                ?           �          �          v       fM     �   �   �   �      6    signal iteration: unsigned(5 downto 0) := "000000"5��    �   6                  M"                     5�_�  *  ,          +   �   .    ����                                                                                                                                                                                                                                                                                                                ?           �          �          v       fP     �   �   �   �      0    counter: counter_6bit port map (clk, rst, );5��    �   .                  �"                     �    �   0                  �"                     �    �   /                  �"                     �    �   .              	   �"             	       �    �   .       	          �"      	              �    �   .              	   �"             	       5�_�  +  M          ,   �       ����                                                                                                                                                                                                                                                                                                                ?           �          �          v       fW     �   �   �   �      7    signal iteration: unsigned(5 downto 0) := "000000";5��    �                    -"                    �    �                     0"                     �    �                     /"                     �    �                     ."                     �    �                    -"                    �    �                     /"                     �    �                     ."                     �    �                 
   -"             
       �    �                     6"                     �    �                     5"                     �    �                     4"                     �    �                     3"                     �    �                     2"                     �    �                     1"                     �    �                     0"                     �    �                     /"                     �    �                     ."                     �    �                 
   -"             
       �    �          
          -"      
              �    �                 
   -"             
       5�_�  ,  N  -      M   =        ����                                                                                                                                                                                                                                                                                                                ?           �          =           V       f�     �   <   =       �           -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );              type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   7        H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   7        H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   7        H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   7        H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   7        H_4 => bit_vector(to_signed(32, 16#510e527f#)),   7        H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   7        H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   6        H_7 => bit_vector(to_signed(32, 16#5be0cd19#))       );5��    <       �               (      �              5�_�  M  O          N   -        ����                                                                                                                                                                                                                                                                                                                            =          =           V       f�     �   ,   �   F    �   -   .   F    5��    ,               �       �              �      5�_�  N  Q          O           ����                                                                                                                                                                                                                                                                                                                            �          �           V       fN     �                use IEEE.STD_LOGIC_1164.ALL;5��                                                5�_�  O  R  P      Q          ����                                                                                                                                                                                                                                                                                                                                                  V        f�     �         �      ,        elsif (clk'event and clk = '1') then5��                        	                    5�_�  Q  S          R          ����                                                                                                                                                                                                                                                                                                                                                  V        f�     �         �              elsif rising_edge then5��                                              5�_�  R  T          S          ����                                                                                                                                                                                                                                                                                                                                                  V        f�    �         �               elsif rising_edge() then5��                                              5�_�  S  U          T   �       ����                                                                                                                                                                                                                                                                                                                                                  V        fm~     �   �   �   �          process�   �   �   �          �   �   �   �    5��    �                      q"                     �    �                      q"                     �    �                     q"                     �    �                     v"                     �    �                     w"                     �    �                    v"                    �    �                    v"                    �    �                    v"                    5�_�  T  V          U   �       ����                                                                                                                                                                                                                                                                                                                                                  V        fm�     �   �   �   �          process5��    �                     }"                     5�_�  U  W          V   �       ����                                                                                                                                                                                                                                                                                                                                                  V        fm�     �   �   �   �          process()5��    �                     ~"                     5�_�  V  X          W   �       ����                                                                                                                                                                                                                                                                                                                                                  V        fm�     �   �   �   �              if rising_edge�   �   �   �          process(clk)5��    �                    �"                     �    �                     �"                    �    �                     �"                    �    �   	                  �"                     �    �   	                  �"                     �    �   	                 �"                     �    �                     �"                    �    �                     �"                     �    �                     �"                     �    �                     �"                     �    �                    �"                    �    �                    �"                    �    �                    �"                    5�_�  W  Y          X   �       ����                                                                                                                                                                                                                                                                                                                                                  V        fm�     �   �   �   �              if rising_edge5��    �                     �"                     5�_�  X  Z          Y   �       ����                                                                                                                                                                                                                                                                                                                                                  V        fm�     �   �   �   �              if rising_edge()5��    �                     �"                     5�_�  Y  [          Z   �       ����                                                                                                                                                                                                                                                                                                                                                  V        fm�     �   �   �   �                  assert�   �   �   �              if rising_edge(clk)5��    �                     �"                     �    �                      �"                     �    �                     �"              	       �    �                     �"                    �    �                     �"                     �    �                     �"                     �    �                    �"                    �    �                    �"                    �    �                    �"                    �    �                 2   �"             2       5�_�  Z  \          [   �       ����                                                                                                                                                                                                                                                                                                                            �          �          v       fm�     �   �   �   �      >            assert neg_condition report message severity note;5��    �                    �"                    5�_�  [  ]          \   �        ����                                                                                                                                                                                                                                                                                                                            �   &       �           v        fm�     �   �   �   �      6            assert false report message severity note;5��    �                     �"                    5�_�  \  ^          ]   �   -    ����                                                                                                                                                                                                                                                                                                                            �   &       �           v        fm�     �   �   �   �      <            assert false report integer'image severity note;5��    �   -                  �"                     5�_�  ]  _          ^   �   .    ����                                                                                                                                                                                                                                                                                                                            �   &       �           v        fm�     �   �   �   �      >            assert false report integer'image() severity note;5��    �   .               
   �"              
       5�_�  ^  `          _   �   8    ����                                                                                                                                                                                                                                                                                                                            �   &       �           v        fm�     �   �   �   �      H            assert false report integer'image(to_integer) severity note;5��    �   8                  �"                     5�_�  _  a          `   �   9    ����                                                                                                                                                                                                                                                                                                                            �   &       �           v        fm�     �   �   �   �      J            assert false report integer'image(to_integer()) severity note;5��    �   9                  �"                     �    �   <                  �"                     �    �   ;                  �"                     �    �   :                  �"                     �    �   9                 �"                    �    �   9                 �"                    �    �   9                 �"                    5�_�  `  b          a   �   A    ����                                                                                                                                                                                                                                                                                                                            �   &       �           v        fm�     �   �   �   �      R            assert false report integer'image(to_integer(unsigned)) severity note;5��    �   A                  �"                     5�_�  a  c          b   �   B    ����                                                                                                                                                                                                                                                                                                                            �   &       �           v        fm�     �   �   �   �      T            assert false report integer'image(to_integer(unsigned())) severity note;5��    �   B                  �"                     �    �   C                  �"                     �    �   B              	   �"             	       �    �   B       	          �"      	              �    �   B              	   �"             	       5�_�  b  d          c   �   I    ����                                                                                                                                                                                                                                                                                                                            �   &       �           v        fm�    �   �   �   �          end process�   �   �   �                  �   �   �   �    5��    �                      #                     �    �                     #                     �    �                    #                    �    �                     #                    �    �                     #                     �    �                    #              	       �    �                     $#                     �    �                     #                    �    �                     $#                     �    �   
                  &#                     �    �   	                  %#                     �    �                    $#                    �    �                    $#                    �    �                    $#                    5�_�  c  e          d   r        ����                                                                                                                                                                                                                                                                                                                /           r          �          V       fnX    �   �   �          6        H_7 => bit_vector(to_signed(32, 16#5be0cd19#))�   �   �          7        H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),�   �   �          7        H_5 => bit_vector(to_signed(32, 16#9b05688c#)),�   �   �          7        H_4 => bit_vector(to_signed(32, 16#510e527f#)),�   �   �          7        H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),�   �   �          7        H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),�   �   �          7        H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),�   �   �          7        H_0 => bit_vector(to_signed(32, 16#6a09e667#)),�   �   �          7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))�   �   �          8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),�   �   �          8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),�   �   �          8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),�   �   �          8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),�   �   �          8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),�   �   �          8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),�   �   �          8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),�   �   �          8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),�   �   �          8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),�   �   �          8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),�   �   �          8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),�   �   �          8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),�   �   �          8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),�   �   �          8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),�   �   �          8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),�   �   �          8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),�   �   �          8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),�   �   �          8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),�   �   �          8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),�   �   �          8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),�   �   �          8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),�   �   �          8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),�   �   �          8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),�   �   �          8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),�   �   �          8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),�   �   �          8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),�   �   �          8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),�   �   �          8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),�   �   �          8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),�   �   �          8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),�   �   �          8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),�   �   �          8        K_31 => bit_vector(to_signed(32, 16#14292967#)),�   �   �          8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),�   �   �          8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),�   �   �          8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),�   �   �          8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),�   �   �          8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),�   �   �          8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),�   �   �          8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),�   �   �          8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),�   �   �          8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),�   �   �          8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),�   �   �          8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),�   �   �          8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),�   �   �          8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),�   �   �          8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),�   �   �          8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),�   �   �          8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),�      �          8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),�   ~   �          8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),�   }             8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),�   |   ~          8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),�   {   }          8        K_10 => bit_vector(to_signed(32, 16#243185be#)),�   z   |          7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),�   y   {          7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),�   x   z          7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),�   w   y          7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),�   v   x          7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),�   u   w          7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),�   t   v          7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),�   s   u          7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),�   r   t          7        K_1 => bit_vector(to_signed(32, 16#71374491#)),�   q   s   �      7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),5��    q                    H                    �    r                    �                    �    s                    �                    �    t                    �                    �    u                    0                    �    v                    j                    �    w                    �                    �    x                    �                    �    y                                        �    z                    R                    �    {                    �                    �    |                    �                    �    }                                        �    ~                    >                    �                        y                    �    �                    �                    �    �                    �                    �    �                    *                    �    �                    e                    �    �                    �                    �    �                    �                    �    �                                        �    �                    Q                    �    �                    �                    �    �                    �                    �    �                                        �    �                    =                    �    �                    x                    �    �                    �                    �    �                    �                    �    �                    )                    �    �                    d                    �    �                    �                    �    �                    �                    �    �                                        �    �                    P                    �    �                    �                    �    �                    �                    �    �                                        �    �                    <                    �    �                    w                    �    �                    �                    �    �                    �                    �    �                    (                    �    �                    c                    �    �                    �                    �    �                    �                    �    �                                        �    �                    O                    �    �                    �                    �    �                    �                    �    �                                         �    �                    ;                    �    �                    v                    �    �                    �                    �    �                    �                    �    �                    '                    �    �                    b                    �    �                    �                    �    �                    �                    �    �                                        �    �                    N                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                                        �    �                    ;                    �    �                    u                    �    �                    �                    �    �                    �                    �    �                    #                     5�_�  d  g          e          ����                                                                                                                                                                                                                                                                                                                /           r          �          V       fnx     �                use IEEE.STD_LOGIC_1164.ALL;5��                          �                     5�_�  e  h  f      g   ,        ����                                                                                                                                                                                                                                                                                                                .                     �          V       fo�     �   ,   /   �          �   ,   .   �    5��    ,                      �                     �    ,                      �                     �    ,                     �                     �    -                      �                     5�_�  g  i          h   -        ����                                                                                                                                                                                                                                                                                                                0                     �          V       fo�     �   ,   /   �       �   -   .   �    5��    ,                      �                     �    ,                 %   �              Q       5�_�  h  j          i   .        ����                                                                                                                                                                                                                                                                                                                1                     �          V       fo�     �   -   /   �      %signal a : int_array := (1, 2, 3, 4);5��    -                      �                     5�_�  i  k          j   .       ����                                                                                                                                                                                                                                                                                                                1                     �          V       fo�     �   -   /   �      )    signal a : int_array := (1, 2, 3, 4);5��    -                                        �    -                                        5�_�  j  l          k   .       ����                                                                                                                                                                                                                                                                                                                1           .          .          v       fo�     �   -   /   �      0    signal k_vector : int_array := (1, 2, 3, 4);5��    -                                          5�_�  k  m          l   -   	    ����                                                                                                                                                                                                                                                                                                                1           .          .          v       fo�     �   ,   .   �      /    type int_array is array(0 to 3) of integer;5��    ,   	       	          �      	              5�_�  l  o          m   -        ����                                                                                                                                                                                                                                                                                                                1           .          .          v       fp     �   ,   .   �      .    type k_vector is array(0 to 3) of integer;5��    ,                      �                     5�_�  m  p  n      o   -   '    ����                                                                                                                                                                                                                                                                                                                1           -   '       -   -       v   -    fp     �   ,   .   �      /    type k_vector is array(0 to 63) of integer;�   -   .   �    5��    ,   '                 �                    5�_�  o  q          p   .       ����                                                                                                                                                                                                                                                                                                                1           -   '       -   =       v   -    fp%     �   -   /   �      )    signal k : int_array := (1, 2, 3, 4);5��    -          	                	              5�_�  p  r          q   .       ����                                                                                                                                                                                                                                                                                                                1           -   '       -   =       v   -    fp.     �   -   0   �      (    signal k : k_vector := (1, 2, 3, 4);5��    -                    (                     5�_�  q  s          r   /       ����                                                                                                                                                                                                                                                                                                                2           -   '       -   =       v   -    fp1     �   .   1   �          1, 2, 3, 4);5��    .                    0                     5�_�  r  t          s   0       ����                                                                                                                                                                                                                                                                                                                3           -   '       -   =       v   -    fp3     �   /   2   �          2, 3, 4);5��    /                    8                     5�_�  s  u          t   1       ����                                                                                                                                                                                                                                                                                                                4           -   '       -   =       v   -    fp6     �   0   3   �      
    3, 4);5��    0                    @                     5�_�  t  v          u   /       ����                                                                                                                                                                                                                                                                                                                5           /          2                 fpP     �   .   4   �                                  ;    �   /   0   �    �   .   3   �          1,        2,        3,        4);5��    .                     -                     �    /                     3                     �    0                     9                     �    1                     ?                     �    .                  *   -              *       �    /                  *   ]              *       �    0                  *   �              *       �    1                  *   �              *       5�_�  u  w          v   2   /    ����                                                                                                                                                                                                                                                                                                                5           /          2   -              fpR     �   1   3   �      /    bit_vector(to_unsigned(32, 16#e9b5dba5#)),;5��    1   .                  �                     �    1   -                 �                    5�_�  v  x          w   2   -    ����                                                                                                                                                                                                                                                                                                                5           /          2   -              fpV     �   1   3   �      .    bit_vector(to_unsigned(32, 16#e9b5dba5#));5��    1   -                  �                     5�_�  w  y          x   2   -    ����                                                                                                                                                                                                                                                                                                                5           /          2   -              fpa     �   1   4   �      /    bit_vector(to_unsigned(32, 16#e9b5dba5#)));5��    1   -                 �                     �    2                      �                     5�_�  x  z          y   3        ����                                                                                                                                                                                                                                                                                                                6           /          2   -              fpc     �   2   4   �      );5��    2                      �                     5�_�  y  |          z   y       ����                                                                                                                                                                                                                                                                                                                6           y          �                 fp}     �   y   �   �   	   9        K_1 => bit_vector(to_unsigned(32, 16#71374491#)),   9        K_2 => bit_vector(to_unsigned(32, 16#b5c0fbcf#)),   9        K_3 => bit_vector(to_unsigned(32, 16#e9b5dba5#)),   9        K_4 => bit_vector(to_unsigned(32, 16#3956c25b#)),   9        K_5 => bit_vector(to_unsigned(32, 16#59f111f1#)),   9        K_6 => bit_vector(to_unsigned(32, 16#923f82a4#)),   9        K_7 => bit_vector(to_unsigned(32, 16#ab1c5ed5#)),   9        K_8 => bit_vector(to_unsigned(32, 16#d807aa98#)),   9        K_9 => bit_vector(to_unsigned(32, 16#12835b01#)),�   x   z   �      9        K_0 => bit_vector(to_unsigned(32, 16#428a2f98#)),5��    x                     @                     �    y                     {                     �    z                     �                     �    {                     �                     �    |                     ,                     �    }                     g                     �    ~                     �                     �                         �                     �    �                                          �    �                     S                     5�_�  z  }  {      |   /       ����                                                                                                                                                                                                                                                                                                                6           2          /   -          -    fp�     �   .   /          /    bit_vector(to_unsigned(32, 16#428a2f98#)),    /    bit_vector(to_unsigned(32, 16#71374491#)), 5��    .                      )      `               5�_�  |            }   /       ����                                                                                                                                                                                                                                                                                                                4           0          /   -          -    fp�     �   .   /          /    bit_vector(to_unsigned(32, 16#b5c0fbcf#)),    -    bit_vector(to_unsigned(32, 16#e9b5dba5#))5��    .                      )      ^               5�_�  }  �  ~         .       ����                                                                                                                                                                                                                                                                                                                2           u          �   9          9    fp�     �   .   0   �    5��    .                      )                     �    .                      )                     5�_�    �  �      �   /        ����                                                                                                                                                                                                                                                                                                                3           v           �           V        fp�     �   /   p   �    �   /   0   �    5��    /               @       *              �      5�_�  �  �          �   /        ����                                                                                                                                                                                                                                                                                                                s           �           �           V        fp�     �   .   /           5��    .                      )                     5�_�  �  �          �   /       ����                                                                                                                                                                                                                                                                                                                r           /          n                 fp�     �   .   o  ,   @   :        K_0 =>  bit_vector(to_unsigned(32, 16#428a2f98#)),   :        K_1 =>  bit_vector(to_unsigned(32, 16#71374491#)),   :        K_2 =>  bit_vector(to_unsigned(32, 16#b5c0fbcf#)),   :        K_3 =>  bit_vector(to_unsigned(32, 16#e9b5dba5#)),   :        K_4 =>  bit_vector(to_unsigned(32, 16#3956c25b#)),   :        K_5 =>  bit_vector(to_unsigned(32, 16#59f111f1#)),   :        K_6 =>  bit_vector(to_unsigned(32, 16#923f82a4#)),   :        K_7 =>  bit_vector(to_unsigned(32, 16#ab1c5ed5#)),   :        K_8 =>  bit_vector(to_unsigned(32, 16#d807aa98#)),   :        K_9 =>  bit_vector(to_unsigned(32, 16#12835b01#)),   :        K_10 => bit_vector(to_unsigned(32, 16#243185be#)),   :        K_11 => bit_vector(to_unsigned(32, 16#550c7dc3#)),   :        K_12 => bit_vector(to_unsigned(32, 16#72be5d74#)),   :        K_13 => bit_vector(to_unsigned(32, 16#80deb1fe#)),   :        K_14 => bit_vector(to_unsigned(32, 16#9bdc06a7#)),   :        K_15 => bit_vector(to_unsigned(32, 16#c19bf174#)),   :        K_16 => bit_vector(to_unsigned(32, 16#e49b69c1#)),   :        K_17 => bit_vector(to_unsigned(32, 16#efbe4786#)),   :        K_18 => bit_vector(to_unsigned(32, 16#0fc19dc6#)),   :        K_19 => bit_vector(to_unsigned(32, 16#240ca1cc#)),   :        K_20 => bit_vector(to_unsigned(32, 16#2de92c6f#)),   :        K_21 => bit_vector(to_unsigned(32, 16#4a7484aa#)),   :        K_22 => bit_vector(to_unsigned(32, 16#5cb0a9dc#)),   :        K_23 => bit_vector(to_unsigned(32, 16#76f988da#)),   :        K_24 => bit_vector(to_unsigned(32, 16#983e5152#)),   :        K_25 => bit_vector(to_unsigned(32, 16#a831c66d#)),   :        K_26 => bit_vector(to_unsigned(32, 16#b00327c8#)),   :        K_27 => bit_vector(to_unsigned(32, 16#bf597fc7#)),   :        K_28 => bit_vector(to_unsigned(32, 16#c6e00bf3#)),   :        K_29 => bit_vector(to_unsigned(32, 16#d5a79147#)),   :        K_30 => bit_vector(to_unsigned(32, 16#06ca6351#)),   :        K_31 => bit_vector(to_unsigned(32, 16#14292967#)),   :        K_32 => bit_vector(to_unsigned(32, 16#27b70a85#)),   :        K_33 => bit_vector(to_unsigned(32, 16#2e1b2138#)),   :        K_34 => bit_vector(to_unsigned(32, 16#4d2c6dfc#)),   :        K_35 => bit_vector(to_unsigned(32, 16#53380d13#)),   :        K_36 => bit_vector(to_unsigned(32, 16#650a7354#)),   :        K_37 => bit_vector(to_unsigned(32, 16#766a0abb#)),   :        K_38 => bit_vector(to_unsigned(32, 16#81c2c92e#)),   :        K_39 => bit_vector(to_unsigned(32, 16#92722c85#)),   :        K_40 => bit_vector(to_unsigned(32, 16#a2bfe8a1#)),   :        K_41 => bit_vector(to_unsigned(32, 16#a81a664b#)),   :        K_42 => bit_vector(to_unsigned(32, 16#c24b8b70#)),   :        K_43 => bit_vector(to_unsigned(32, 16#c76c51a3#)),   :        K_44 => bit_vector(to_unsigned(32, 16#d192e819#)),   :        K_45 => bit_vector(to_unsigned(32, 16#d6990624#)),   :        K_46 => bit_vector(to_unsigned(32, 16#f40e3585#)),   :        K_47 => bit_vector(to_unsigned(32, 16#106aa070#)),   :        K_48 => bit_vector(to_unsigned(32, 16#19a4c116#)),   :        K_49 => bit_vector(to_unsigned(32, 16#1e376c08#)),   :        K_50 => bit_vector(to_unsigned(32, 16#2748774c#)),   :        K_51 => bit_vector(to_unsigned(32, 16#34b0bcb5#)),   :        K_52 => bit_vector(to_unsigned(32, 16#391c0cb3#)),   :        K_53 => bit_vector(to_unsigned(32, 16#4ed8aa4a#)),   :        K_54 => bit_vector(to_unsigned(32, 16#5b9cca4f#)),   :        K_55 => bit_vector(to_unsigned(32, 16#682e6ff3#)),   :        K_56 => bit_vector(to_unsigned(32, 16#748f82ee#)),   :        K_57 => bit_vector(to_unsigned(32, 16#78a5636f#)),   :        K_58 => bit_vector(to_unsigned(32, 16#84c87814#)),   :        K_59 => bit_vector(to_unsigned(32, 16#8cc70208#)),   :        K_60 => bit_vector(to_unsigned(32, 16#90befffa#)),   :        K_61 => bit_vector(to_unsigned(32, 16#a4506ceb#)),   :        K_62 => bit_vector(to_unsigned(32, 16#bef9a3f7#)),   9        K_63 => bit_vector(to_unsigned(32, 16#c67178f2#))5��    .                     1                     �    /                     d                     �    0                     �                     �    1                     �                     �    2                     �                     �    3                     0                     �    4                     c                     �    5                     �                     �    6                     �                     �    7                     �                     �    8                     /                     �    9                     b                     �    :                     �                     �    ;                     �                     �    <                     �                     �    =                     .                     �    >                     a                     �    ?                     �                     �    @                     �                     �    A                     �                     �    B                     -                     �    C                     `                     �    D                     �                     �    E                     �                     �    F                     �                     �    G                     ,	                     �    H                     _	                     �    I                     �	                     �    J                     �	                     �    K                     �	                     �    L                     +
                     �    M                     ^
                     �    N                     �
                     �    O                     �
                     �    P                     �
                     �    Q                     *                     �    R                     ]                     �    S                     �                     �    T                     �                     �    U                     �                     �    V                     )                     �    W                     \                     �    X                     �                     �    Y                     �                     �    Z                     �                     �    [                     (                     �    \                     [                     �    ]                     �                     �    ^                     �                     �    _                     �                     �    `                     '                     �    a                     Z                     �    b                     �                     �    c                     �                     �    d                     �                     �    e                     &                     �    f                     Y                     �    g                     �                     �    h                     �                     �    i                     �                     �    j                     %                     �    k                     X                     �    l                     �                     �    m                     �                     5�_�  �  �          �   q        ����                                                                                                                                                                                                                                                                                                                r           q          �          V       fp�     �   p   q       �       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   :        K_0 =>  bit_vector(to_unsigned(32, 16#428a2f98#)),   :        K_1 =>  bit_vector(to_unsigned(32, 16#71374491#)),   :        K_2 =>  bit_vector(to_unsigned(32, 16#b5c0fbcf#)),   :        K_3 =>  bit_vector(to_unsigned(32, 16#e9b5dba5#)),   :        K_4 =>  bit_vector(to_unsigned(32, 16#3956c25b#)),   :        K_5 =>  bit_vector(to_unsigned(32, 16#59f111f1#)),   :        K_6 =>  bit_vector(to_unsigned(32, 16#923f82a4#)),   :        K_7 =>  bit_vector(to_unsigned(32, 16#ab1c5ed5#)),   :        K_8 =>  bit_vector(to_unsigned(32, 16#d807aa98#)),   :        K_9 =>  bit_vector(to_unsigned(32, 16#12835b01#)),   :        K_10 => bit_vector(to_unsigned(32, 16#243185be#)),   :        K_11 => bit_vector(to_unsigned(32, 16#550c7dc3#)),   :        K_12 => bit_vector(to_unsigned(32, 16#72be5d74#)),   :        K_13 => bit_vector(to_unsigned(32, 16#80deb1fe#)),   :        K_14 => bit_vector(to_unsigned(32, 16#9bdc06a7#)),   :        K_15 => bit_vector(to_unsigned(32, 16#c19bf174#)),   :        K_16 => bit_vector(to_unsigned(32, 16#e49b69c1#)),   :        K_17 => bit_vector(to_unsigned(32, 16#efbe4786#)),   :        K_18 => bit_vector(to_unsigned(32, 16#0fc19dc6#)),   :        K_19 => bit_vector(to_unsigned(32, 16#240ca1cc#)),   :        K_20 => bit_vector(to_unsigned(32, 16#2de92c6f#)),   :        K_21 => bit_vector(to_unsigned(32, 16#4a7484aa#)),   :        K_22 => bit_vector(to_unsigned(32, 16#5cb0a9dc#)),   :        K_23 => bit_vector(to_unsigned(32, 16#76f988da#)),   :        K_24 => bit_vector(to_unsigned(32, 16#983e5152#)),   :        K_25 => bit_vector(to_unsigned(32, 16#a831c66d#)),   :        K_26 => bit_vector(to_unsigned(32, 16#b00327c8#)),   :        K_27 => bit_vector(to_unsigned(32, 16#bf597fc7#)),   :        K_28 => bit_vector(to_unsigned(32, 16#c6e00bf3#)),   :        K_29 => bit_vector(to_unsigned(32, 16#d5a79147#)),   :        K_30 => bit_vector(to_unsigned(32, 16#06ca6351#)),   :        K_31 => bit_vector(to_unsigned(32, 16#14292967#)),   :        K_32 => bit_vector(to_unsigned(32, 16#27b70a85#)),   :        K_33 => bit_vector(to_unsigned(32, 16#2e1b2138#)),   :        K_34 => bit_vector(to_unsigned(32, 16#4d2c6dfc#)),   :        K_35 => bit_vector(to_unsigned(32, 16#53380d13#)),   :        K_36 => bit_vector(to_unsigned(32, 16#650a7354#)),   :        K_37 => bit_vector(to_unsigned(32, 16#766a0abb#)),   :        K_38 => bit_vector(to_unsigned(32, 16#81c2c92e#)),   :        K_39 => bit_vector(to_unsigned(32, 16#92722c85#)),   :        K_40 => bit_vector(to_unsigned(32, 16#a2bfe8a1#)),   :        K_41 => bit_vector(to_unsigned(32, 16#a81a664b#)),   :        K_42 => bit_vector(to_unsigned(32, 16#c24b8b70#)),   :        K_43 => bit_vector(to_unsigned(32, 16#c76c51a3#)),   :        K_44 => bit_vector(to_unsigned(32, 16#d192e819#)),   :        K_45 => bit_vector(to_unsigned(32, 16#d6990624#)),   :        K_46 => bit_vector(to_unsigned(32, 16#f40e3585#)),   :        K_47 => bit_vector(to_unsigned(32, 16#106aa070#)),   :        K_48 => bit_vector(to_unsigned(32, 16#19a4c116#)),   :        K_49 => bit_vector(to_unsigned(32, 16#1e376c08#)),   :        K_50 => bit_vector(to_unsigned(32, 16#2748774c#)),   :        K_51 => bit_vector(to_unsigned(32, 16#34b0bcb5#)),   :        K_52 => bit_vector(to_unsigned(32, 16#391c0cb3#)),   :        K_53 => bit_vector(to_unsigned(32, 16#4ed8aa4a#)),   :        K_54 => bit_vector(to_unsigned(32, 16#5b9cca4f#)),   :        K_55 => bit_vector(to_unsigned(32, 16#682e6ff3#)),   :        K_56 => bit_vector(to_unsigned(32, 16#748f82ee#)),   :        K_57 => bit_vector(to_unsigned(32, 16#78a5636f#)),   :        K_58 => bit_vector(to_unsigned(32, 16#84c87814#)),   :        K_59 => bit_vector(to_unsigned(32, 16#8cc70208#)),   :        K_60 => bit_vector(to_unsigned(32, 16#90befffa#)),   :        K_61 => bit_vector(to_unsigned(32, 16#a4506ceb#)),   :        K_62 => bit_vector(to_unsigned(32, 16#bef9a3f7#)),   9        K_63 => bit_vector(to_unsigned(32, 16#c67178f2#))       );5��    p       �               �                    5�_�  �  �          �   q       ����                                                                                                                                                                                                                                                                                                                            q          q          V       fp�    �   p   q              5��    p                      �                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       fq    �   �   �   �          process(clk)   	    begin            if rising_edge(clk) then   ]            assert false report integer'image(to_integer(unsigned(iteration))) severity note;           end if;       end process;5��    �                           �       �       5�_�  �  �  �      �   ,       ����                                                                                                                                                                                                                                                                                                                            �          ,          V   -    fr�     �   +   ,       Z       -- Constants   ?    type k_vector is array(0 to 63) of bit_vector(31 downto 0);       signal k : k_vector := (   2        bit_vector(to_unsigned(32, 16#428a2f98#)),   2        bit_vector(to_unsigned(32, 16#71374491#)),   2        bit_vector(to_unsigned(32, 16#b5c0fbcf#)),   2        bit_vector(to_unsigned(32, 16#e9b5dba5#)),   2        bit_vector(to_unsigned(32, 16#3956c25b#)),   2        bit_vector(to_unsigned(32, 16#59f111f1#)),   2        bit_vector(to_unsigned(32, 16#923f82a4#)),   2        bit_vector(to_unsigned(32, 16#ab1c5ed5#)),   2        bit_vector(to_unsigned(32, 16#d807aa98#)),   2        bit_vector(to_unsigned(32, 16#12835b01#)),   2        bit_vector(to_unsigned(32, 16#243185be#)),   2        bit_vector(to_unsigned(32, 16#550c7dc3#)),   2        bit_vector(to_unsigned(32, 16#72be5d74#)),   2        bit_vector(to_unsigned(32, 16#80deb1fe#)),   2        bit_vector(to_unsigned(32, 16#9bdc06a7#)),   2        bit_vector(to_unsigned(32, 16#c19bf174#)),   2        bit_vector(to_unsigned(32, 16#e49b69c1#)),   2        bit_vector(to_unsigned(32, 16#efbe4786#)),   2        bit_vector(to_unsigned(32, 16#0fc19dc6#)),   2        bit_vector(to_unsigned(32, 16#240ca1cc#)),   2        bit_vector(to_unsigned(32, 16#2de92c6f#)),   2        bit_vector(to_unsigned(32, 16#4a7484aa#)),   2        bit_vector(to_unsigned(32, 16#5cb0a9dc#)),   2        bit_vector(to_unsigned(32, 16#76f988da#)),   2        bit_vector(to_unsigned(32, 16#983e5152#)),   2        bit_vector(to_unsigned(32, 16#a831c66d#)),   2        bit_vector(to_unsigned(32, 16#b00327c8#)),   2        bit_vector(to_unsigned(32, 16#bf597fc7#)),   2        bit_vector(to_unsigned(32, 16#c6e00bf3#)),   2        bit_vector(to_unsigned(32, 16#d5a79147#)),   2        bit_vector(to_unsigned(32, 16#06ca6351#)),   2        bit_vector(to_unsigned(32, 16#14292967#)),   2        bit_vector(to_unsigned(32, 16#27b70a85#)),   2        bit_vector(to_unsigned(32, 16#2e1b2138#)),   2        bit_vector(to_unsigned(32, 16#4d2c6dfc#)),   2        bit_vector(to_unsigned(32, 16#53380d13#)),   2        bit_vector(to_unsigned(32, 16#650a7354#)),   2        bit_vector(to_unsigned(32, 16#766a0abb#)),   2        bit_vector(to_unsigned(32, 16#81c2c92e#)),   2        bit_vector(to_unsigned(32, 16#92722c85#)),   2        bit_vector(to_unsigned(32, 16#a2bfe8a1#)),   2        bit_vector(to_unsigned(32, 16#a81a664b#)),   2        bit_vector(to_unsigned(32, 16#c24b8b70#)),   2        bit_vector(to_unsigned(32, 16#c76c51a3#)),   2        bit_vector(to_unsigned(32, 16#d192e819#)),   2        bit_vector(to_unsigned(32, 16#d6990624#)),   2        bit_vector(to_unsigned(32, 16#f40e3585#)),   2        bit_vector(to_unsigned(32, 16#106aa070#)),   2        bit_vector(to_unsigned(32, 16#19a4c116#)),   2        bit_vector(to_unsigned(32, 16#1e376c08#)),   2        bit_vector(to_unsigned(32, 16#2748774c#)),   2        bit_vector(to_unsigned(32, 16#34b0bcb5#)),   2        bit_vector(to_unsigned(32, 16#391c0cb3#)),   2        bit_vector(to_unsigned(32, 16#4ed8aa4a#)),   2        bit_vector(to_unsigned(32, 16#5b9cca4f#)),   2        bit_vector(to_unsigned(32, 16#682e6ff3#)),   2        bit_vector(to_unsigned(32, 16#748f82ee#)),   2        bit_vector(to_unsigned(32, 16#78a5636f#)),   2        bit_vector(to_unsigned(32, 16#84c87814#)),   2        bit_vector(to_unsigned(32, 16#8cc70208#)),   2        bit_vector(to_unsigned(32, 16#90befffa#)),   2        bit_vector(to_unsigned(32, 16#a4506ceb#)),   2        bit_vector(to_unsigned(32, 16#bef9a3f7#)),   1        bit_vector(to_unsigned(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   9        H_0 => bit_vector(to_unsigned(32, 16#6a09e667#)),   9        H_1 => bit_vector(to_unsigned(32, 16#bb67ae85#)),   9        H_2 => bit_vector(to_unsigned(32, 16#3c6ef372#)),   9        H_3 => bit_vector(to_unsigned(32, 16#a54ff53a#)),   9        H_4 => bit_vector(to_unsigned(32, 16#510e527f#)),   9        H_5 => bit_vector(to_unsigned(32, 16#9b05688c#)),   9        H_6 => bit_vector(to_unsigned(32, 16#1f83d9ab#)),   8        H_7 => bit_vector(to_unsigned(32, 16#5be0cd19#))       );5��    +       Z               �      �              5�_�  �  �          �   ,        ����                                                                                                                                                                                                                                                                                                                            ,          ,          V   -    fr�    �   +   ,           5��    +                      �                     5�_�  �  �          �   C        ����                                                                                                                                                                                                                                                                                                                            H           C           V        fr�    �   B   I   K          -- process(clk)       -- begin   #    --     if rising_edge(clk) then   `    --         assert false report integer'image(to_integer(unsigned(iteration))) severity note;       --     end if;       -- end process;5��    B                     v      �       �       5�_�  �  �          �   =        ����                                                                                                                                                                                                                                                                                                                            H           C           V        fs     �   =   ?   K    �   =   >   K    5��    =                      /              .       5�_�  �  �          �   >       ����                                                                                                                                                                                                                                                                                                                            I           D           V        fs     �   =   ?   L      -    signal clk : bit := '0';  -- Clock signal5��    =                    :                    5�_�  �  �          �   B   $    ����                                                                                                                                                                                                                                                                                                                            I           D           V        fs     �   A   C   L      9    counter: counter_6bit port map (clk, rst, iteration);5��    A   $                 �                    5�_�  �  �          �   D       ����                                                                                                                                                                                                                                                                                                                            I           D           V        fs     �   C   E   L          process(clk)5��    C                    �                    5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                            I           D           V        fs     �   E   G   L               if rising_edge(clk) then5��    E                    �                    5�_�  �  �          �   @       ����                                                                                                                                                                                                                                                                                                                            I           D           V        fs%     �   @   K   L    �   @   A   L    5��    @               
       f              �       5�_�  �  �          �   D       ����                                                                                                                                                                                                                                                                                                                            S           N           V        fs(     �   C   E   V              clk <= '0';5��    C                    �                    5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            S           N           V        fs.     �   F   H   V                  clk <= not clk;5��    F                    �                    5�_�  �  �          �   ;        ����                                                                                                                                                                                                                                                                                                                            S           N           V        fs>    �   ;   =   V    �   ;   <   V    5��    ;                      �              K       5�_�  �  �          �   Q       ����                                                                                                                                                                                                                                                                                                                            T           O           V        fu     �   Q   S   W    �   Q   R   W    5��    Q                      0              '       5�_�  �  �  �      �   R       ����                                                                                                                                                                                                                                                                                                                            U           O           V        fuv     �   Q   R          &            wait for CLOCK_PERIOD / 2;5��    Q                      0      '               5�_�  �  �          �   Q       ����                                                                                                                                                                                                                                                                                                                            T           O           V        fuw     �   P   R   X              �   P   R   W    5��    P                                    	       �    P                                          �    P                 	                	       5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                            R          T                 fu�     �   R   U   X      ]            assert false report integer'image(to_integer(unsigned(iteration))) severity note;           end if;�   Q   S   X      "        if rising_edge(clock) then5��    Q                     -                     �    R                     T                     �    S                     �                     5�_�  �  �          �   T       ����                                                                                                                                                                                                                                                                                                                            R          T                 fu�    �   T   V   Y                  �   T   V   X    5��    T                      �                     �    T                     �                     �    T                     �                    �    T                     �                     5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                            R          T                 fu�     �   Q   R          &            if rising_edge(clock) then5��    Q                      %      '               5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                            R          S                 fu�     �   R   S                      end if;5��    R                      �                     5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                            R          S                 fu�    �   Q   S   W      a                assert false report integer'image(to_integer(unsigned(iteration))) severity note;5��    Q                     1                     5�_�  �  �  �      �   <        ����                                                                                                                                                                                                                                                                                                                            #          &          V       f��     �   ;   <          J    constant CLOCK_PERIOD : time := 20 ns;  -- Clock period (e.g., 50 MHz)5��    ;                      �      K               5�_�  �  �          �   >        ����                                                                                                                                                                                                                                                                                                                            #          &          V       f��     �   =   >          /    signal clock : bit := '0';  -- Clock signal5��    =                      /      0               5�_�  �  �          �   @        ����                                                                                                                                                                                                                                                                                                                            @           I           V        f��     �   ?   @       
       -- Clock process       clk_process: process   	    begin           clock <= '0';   "        wait for CLOCK_PERIOD / 2;           while true loop               clock <= not clk;   &            wait for CLOCK_PERIOD / 2;           end loop;       end process clk_process;5��    ?       
               6      �               5�_�  �  �          �   A   $    ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��     �   @   B   K      ;    counter: counter_6bit port map (clock, rst, iteration);5��    @   $                 _                    5�_�  �  �          �   C       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��    �   B   D   K          process(clock)5��    B                    �                    �    B                    �                    5�_�  �  �  �      �   E       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f�	     �   D   E                  while true loop5��    D                      �                     5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f�     �   E   F                  end loop;5��    E                      �                     5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f�    �   D   F   I      ]            assert false report integer'image(to_integer(unsigned(iteration))) severity note;5��    D                     �                     5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��     �   D   F   I      Y        assert false report integer'image(to_integer(unsigned(iteration))) severity note;5��    D                    �                    �    D                     �                     �    D                 	   �             	       �    D          	          �      	              �    D                    �                    5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��     �   D   F   I      `        assert iteration =  report integer'image(to_integer(unsigned(iteration))) severity note;5��    D                     �                     5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��     �   D   F   I      b        assert iteration = "" report integer'image(to_integer(unsigned(iteration))) severity note;5��    D                     �                     5�_�  �  �          �   E        ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��     �   D   F   I      h        assert iteration = "000000" report integer'image(to_integer(unsigned(iteration))) severity note;5��    D                     �                    5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��     �   D   F   I      h        assert iteration = "000010" report integer'image(to_integer(unsigned(iteration))) severity note;5��    D                     �                     5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��   ! �   D   F   I      i        assert iteration != "000010" report integer'image(to_integer(unsigned(iteration))) severity note;5��    D                    �                    5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��     �   F   H   K              if iteration�   E   H   J              �   E   G   I    5��    E                      �              	       �    E                      �                     �    E                     �              	       �    F                                          �    F                                          �    F                 	                	       �    F          	                	              �    F                                        5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��     �   F   H   K              if iteration = 5��    F                                          5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��     �   F   H   K              if iteration = ""5��    F                                          5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��     �   F   I   K              if iteration = "000000"5��    F                                          �    F                                         �    F   $                                        �    F   $                                	       �    G                     !                    �    G                     -                     5�_�  �  �          �   =       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f�I     �   =   ?   M          �   =   ?   L    5��    =                      /                     �    =                  	   3              	       �    =                    ;                    �    =                    ;                    �    =                     ?                     �    =                     >                     �    =                    =                    �    =                     ?                     �    =                     >                     �    =                 
   =             
       �    =                     F                     �    =                     E                     �    =                     D                     �    =                     C                     �    =                     B                     �    =                     A                     �    =                     @                     �    =                     ?                     �    =                     >                     �    =                 
   =             
       �    =          
          =      
              �    =                 
   =             
       5�_�  �  �          �   >       ����                                                                                                                                                                                                                                                                                                                            A           A           V        f�X     �   =   ?   M          signal w: bit_vector5��    =                     G                     5�_�  �  �          �   >       ����                                                                                                                                                                                                                                                                                                                            A           A           V        f�d     �   =   ?   M          signal w: bit_vector()5��    =                     H                     �    =                    L                    �    =                    L                    �    =                    L                    5�_�  �  �          �   >   &    ����                                                                                                                                                                                                                                                                                                                            A           A           V        f�i     �   =   ?   M      &    signal w: bit_vector(511 downto 0)5��    =   &                  U                     �    =   +                  Z                     �    =   *                 Y                    �    =   *                 Y                    �    =   *                 Y                    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            A           A           V        f�     �      	   M      Q        count : out bit_vector(5 downto 0)       -- 6-bit count output (64 steps)5��                        �                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            A           A           V        f�     �         M      !    count <= bit_vector(counter);5��              
       
   l      
       
       5�_�  �  �          �   8       ����                                                                                                                                                                                                                                                                                                                            A           A           V        f�|     �   7   9   M      U            count : out bit_vector(5 downto 0)       -- 6-bit count output (64 steps)5��    7                    z                    5�_�  �  �          �   =   /    ����                                                                                                                                                                                                                                                                                                                            A           A           V        f��     �   <   >   M      9    signal iteration: bit_vector(5 downto 0) := "000000";5��    <   /       	                	              5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                            A           A           V        f��     �   E   G   M      i        assert iteration /= "000010" report integer'image(to_integer(unsigned(iteration))) severity note;5��    E          	          �      	              5�_�  �  �          �   H       ����                                                                                                                                                                                                                                                                                                                            A           A           V        f��     �   G   H          $        if iteration = "000000" then5��    G                             %               5�_�  �  �          �   H       ����                                                                                                                                                                                                                                                                                                                            A           A           V        f��     �   G   H                      5��    G                                            5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                            A           A           V        f��     �   E   G   K      b        assert iteration /= 2 report integer'image(to_integer(unsigned(iteration))) severity note;5��    E                    �                    5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                            A           A           V        f��     �   E   G   K      b        assert iteration != 2 report integer'image(to_integer(unsigned(iteration))) severity note;5��    E                     �                     5�_�  �  �          �   =       ����                                                                                                                                                                                                                                                                                                                            A           A           V        f��     �   <   >   K      2    signal iteration: bit_vector(5 downto 0) := 0;5��    <                    �                    5�_�  �  �          �   F   2    ����                                                                                                                                                                                                                                                                                                                            A           A           V        f��   " �   E   G   K      a        assert iteration = 2 report integer'image(to_integer(unsigned(iteration))) severity note;5��    E   2                 �                    �    E   3                  �                     �    E   2              	   �             	       �    E   2       	          �      	              �    E   2              	   �             	       5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f��     �   G   J   M              if iteration�   F   I   L              �   F   H   K    5��    F                      �              	       �    F                      �                     �    F                     �              	       �    G                     �                     �    G                     �                     �    G                 	   �             	       �    G          	          �      	              �    G                    �                    �    G                    �                    �    G                    �                    �    G                    �                    �    G                    �              	       �    H                     �                    �    H                     �                    �    H                                          �    H                     �                    �    H                                          5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f��     �   H   J   N                  end if;5��    H                                          5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f��     �   E   F          K        assert iteration = 2 report integer'image(iteration) severity note;5��    E                      �      L               5�_�  �  �          �   G        ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f��     �   G   I   M    �   G   H   M    5��    G                      �              L       5�_�  �  �          �   H       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f��     �   G   I   N      K        assert iteration = 2 report integer'image(iteration) severity note;5��    G                     �                     5�_�  �  �          �   H       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f��   # �   G   I   N      O            assert iteration = 2 report integer'image(iteration) severity note;5��    G                    �                    5�_�  �  �          �   >       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�#     �   =   ?   N      /    signal w: bit_vector(511 downto 0) := msgi;5��    =                                          5�_�  �  �          �   >       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�&     �   >   @   O          �   >   @   N    5��    >                      2                     �    >                     6                     �    >                     B                     �    >                     A                     �    >                    @                    �    >                     B                     �    >                     A                     �    >                 
   @             
       �    >                     I                     �    >                     H                     �    >                     G                     �    >                     F                     �    >                     E                     �    >                     D                     �    >                     C                     �    >                     B                     �    >                     A                     �    >                 
   @             
       �    >          
          @      
              �    >                 
   @             
       5�_�  �  �          �   ?       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�7     �   >   @   O          signal w: bit_vector5��    >                     J                     5�_�  �  �          �   ?       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�:     �   >   @   O          signal w: bit_vector()5��    >                     K                     �    >                    N                    �    >                    N                    �    >                    N                    5�_�  �  �          �   ?   %    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�>     �   >   @   O      %    signal w: bit_vector(31 downto 0)5��    >   %                  W                     5�_�  �  �          �   I   %    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f��     �   H   J   P                  �   H   J   O    5��    H                      �                     �    H                  	   �              	       5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f��     �   H   J   P                  w <= msgi5��    H                     �                     5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f��     �   H   J   P                  w <= msgi()5��    H                     �                     �    H                     �                     5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f��     �   H   J   P                  w <= msgi()5��    H                     �                     �    H                    �                    �    H                    �                    �    H                    �                    �    H                    �                    �    H                    �                    5�_�  �  �          �   I   %    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�     �   H   J   P      %            w <= msgi(16 +2 downto 0)5��    H   %                                        5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�     �   H   J   P      &            w <= msgi(16 +2 downto 0);5��    H                    �                    5�_�  �  �          �   I   "    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�     �   H   J   P      %            w <= msgi(16*2 downto 0);5��    H   "                  �                     �    H   #                 �                    5�_�  �  �          �   I   %    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�$     �   H   J   P      '            w <= msgi(16*2 downto i*0);5��    H   $                 �                    5�_�  �  �          �   I   #    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�*     �   H   J   P      (            w <= msgi(16*2 downto i*16);5��    H   #                  �                     �    H   $                  �                     �    H   #                  �                     �    H   "              	   �             	       �    H   "       	          �      	              �    H   "              	   �             	       5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�-     �   H   J   P      0            w <= msgi(16*2 downto iteration*16);5��    H                     �                     5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�0     �   H   J   P      .            w <= msgi(16 downto iteration*16);5��    H                     �                     �    H                     �                     �    H                 	   �             	       �    H          	          �      	              �    H                 
   �             
       5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�6     �   H   J   P      8            w <= msgi(iteration*16 downto iteration*16);5��    H                     �                     5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�9     �   H   J   P      9            w <= msgi((iteration*16 downto iteration*16);5��    H                     �      :       ;       5�_�  �  �          �   I   $    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�=     �   H   J   P      :            w <= msgi((iteration*16) downto iteration*16);5��    H   $                  �                     5�_�  �  �          �   J   .    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�B     �   I   K   P      G            assert false report integer'image(iteration) severity note;5��    I   .       	          F      	              �    I   /                  G                     �    I   .              
   F             
       �    I   .       
          F      
              �    I   .              
   F             
       5�_�  �  �          �   J   8    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�U     �   I   K   P      H            assert false report integer'image(to_integer) severity note;5��    I   8                  P                     5�_�  �  �          �   J   9    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       f�V     �   I   K   P      J            assert false report integer'image(to_integer()) severity note;5��    I   9                  Q                     �    I   :                  R                     �    I   9                 Q                    �    I   9                 Q                    �    I   9                 Q                    �    I   9                 Q                    5�_�  �  �          �   J   B    ����                                                                                                                                                                                                                                                                                                                            J   B       J   B       v   B    f�Z   $ �   I   K   P      ^            assert false report integer'image(to_integer(unsigned(7 downto 0))) severity note;5��    I   B       
          Z      
              5�_�  �  �          �   I   &    ����                                                                                                                                                                                                                                                                                                                            J   B       J   B       v   B    f��   % �   H   J   P      <            w <= msgi((iteration*16)-1 downto iteration*16);5��    H   %                                        �    H   $                 �                    5�_�  �  �  �      �   J   #    ����                                                                                                                                                                                                                                                                                                                            J   B       J   B       v   B    f��     �   J   L   P    �   J   K   P    5��    J                      o              V       5�_�  �  �          �   K       ����                                                                                                                                                                                                                                                                                                                            J   B       J   B       v   B    f��     �   K   M   Q    �   K   L   Q    5��    K                      �              V       5�_�  �  �          �   K   .    ����                                                                                                                                                                                                                                                                                                                            J   B       J   B       v   B    f�      �   J   L   R      U            assert false report integer'image(to_integer(unsigned(w))) severity note;5��    J   .                 �                    �    J   /                  �                     �    J   .              	   �             	       �    J   .       	          �      	              �    J   .                 �                    �    J   9                 �                    �    J   ;                  �                     5�_�  �  �          �   K   .    ����                                                                                                                                                                                                                                                                                                                            J   B       J   B       v   B    f�     �   J   L   R      K            assert false report integer'image(iteration*16)) severity note;5��    J   .                  �                     5�_�  �  �          �   K   <    ����                                                                                                                                                                                                                                                                                                                            J   B       J   B       v   B    f�     �   J   L   R      L            assert false report integer'image((iteration*16)) severity note;5��    J   <                  �                     5�_�  �  �          �   L   .    ����                                                                                                                                                                                                                                                                                                                            J   B       J   B       v   B    f�     �   K   M   R      U            assert false report integer'image(to_integer(unsigned(w))) severity note;5��    K   .                 �                    �    K   /                  �                     �    K   .              	   �             	       �    K   .       	          �      	              �    K   .                 �                    5�_�  �  �          �   L   ;    ����                                                                                                                                                                                                                                                                                                                            J   B       J   B       v   B    f�#     �   K   M   R      L            assert false report integer'image(iteration/1==*) severity note;5��    K   :                  �                     �    K   9                  �                     �    K   8                  �                     �    K   7                  �                     5�_�  �  �          �   L   8    ����                                                                                                                                                                                                                                                                                                                            J   B       J   B       v   B    f�*   & �   K   M   R      H            assert false report integer'image(iteration*) severity note;5��    K   8                  �                     5�_�  �  �  �      �   L   9    ����                                                                                                                                                                                                                                                                                                                            K   9       L   9       V   9    f�R     �   J   M   R      N            assert false report integer'image((iteration*16)+1) severity note;   J            assert false report integer'image(iteration*16) severity note;5��    J                     o      �       �       5�_�  �  �          �   I   9    ����                                                                                                                                                                                                                                                                                                                            K   9       L   9       V   9    f�T   ) �   H   J   R      =            w <= msgi((iteration*16)+15 downto iteration*16);5��    H                     �      >       A       5�_�  �  �          �   I   9    ����                                                                                                                                                                                                                                                                                                                            K   9       L   9       V   9    f�\     �   H   J   R      @            -- w <= msgi((iteration*16)+15 downto iteration*16);5��    H                     �      A       >       5�_�  �  �          �   K   9    ����                                                                                                                                                                                                                                                                                                                            L   9       K   9       V   9    f�`     �   J   M   R      Q            -- assert false report integer'image((iteration*16)+1) severity note;   M            -- assert false report integer'image(iteration*16) severity note;5��    J                     o      �       �       5�_�  �  �          �   K   >    ����                                                                                                                                                                                                                                                                                                                            L   9       K   9       V   9    f�q     �   J   L   R      N            assert false report integer'image((iteration*16)+1) severity note;5��    J   >                  �                     5�_�  �  �          �   J   >    ����                                                                                                                                                                                                                                                                                                                            I   <       J   >       V   >    f��     �   H   K   R      =            w <= msgi((iteration*16)+15 downto iteration*16);   U            assert false report integer'image(to_integer(unsigned(w))) severity note;5��    H                     �      �       �       5�_�  �             �   K   >    ����                                                                                                                                                                                                                                                                                                                            I   <       J   >       V   >    f��   * �   J   L   R      O            assert false report integer'image((iteration*16)+15) severity note;5��    J                     u      P       S       5�_�  �    �          L   8    ����                                                                                                                                                                                                                                                                                                                            L   I       <           v        f��   + �   K   M   R      J            assert false report integer'image(iteration*16) severity note;5��    K   8                                      5�_�                  L   9    ����                                                                                                                                                                                                                                                                                                                            L   I       <           v        f��   , �   K   M   R      I            assert false report integer'image(iteration*2) severity note;5��    K   8                                        �    K   7                 �                    5�_�                 L   9    ����                                                                                                                                                                                                                                                                                                                            L   I       <           v        f�1   - �   K   M   R      I            assert false report integer'image(iteration+2) severity note;5��    K   8                                      5�_�                 =   "    ����                                                                                                                                                                                                                                                                                                                            L   I       <           v        f��     �   <   >   R      #    signal iteration: integer := 0;5��    <   "                  �                     5�_�                 =   "    ����                                                                                                                                                                                                                                                                                                                            =   "       =   3       v   3    f��     �   <   >   R      5    signal iteration: integer := 0 range -512 to 511;5��    <   "                  �                     5�_�                      ����                                                                                                                                                                                                                                                                                                                            =          =          v       f�     �   !   #   U      use IEEE.numeric_std.all;�      #   S       �      !   R    5��                          �                     �                          �                     �                         �                     �                         �                    �                         �                     �                         �                     �                         �                    �                         �                     �                         �                     �                         �                    �                         �                     �                         �                     �                         �                     �                         �                    �                         �                    �                         �                    �                          �                     �                         �              D       �    !                      	                      5�_�                 !       ����                                                                                                                                                                                                                                                                                                                            @          @          v       f�     �       !          use IEEE.std_logic_1164.all;5��                           �                     5�_�    	                     ����                                                                                                                                                                                                                                                                                                                            ?          ?          v       f�     �                 library IEEE;5��                          �                     5�_�    
          	       	    ����                                                                                                                                                                                                                                                                                                                            >          >          v       f�     �      !   S      use IEEE.numeric_std.all;5��       	                 �                    �       
                  �                     �       	                 �                    �                         �                     �                         �                     �       
                  �                     �       	                 �                    �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �       
                  �                     �       	                 �                    �       	                 �                    �       	                 �                    �       	                 �                    5�_�  	            
       	    ����                                                                                                                                                                                                                                                                                                                            >          >          v       f�     �      !   S      use IEEE.std_logic_arith.all;5��       	                 �                    5�_�  
                 
    ����                                                                                                                                                                                                                                                                                                                            >          >          v       f�v     �                 use IEEE.ar.all;5��                          �                     5�_�               L   7    ����                                                                                                                                                                                                                                                                                                                            =          =          v       f��   1 �   K   M   R      K            assert false report integer'image(iteration+800) severity note;5��    K   7                 �                    5�_�                 ?   %    ����                                                                                                                                                                                                                                                                                                                            =          =          v       f��     �   ?   B   S          �   ?   A   R    5��    ?                      Y                     �    ?                      Y                     �    ?                     Y                     �    @                     ^                     �    @                     j                     �    @                     i                     �    @                     h                     �    @                    g                    5�_�                 N   .    ����                                                                                                                                                                                                                                                                                                                            =          =          v       f�   2 �   M   O   T      I            assert false report integer'image(iteration*2) severity note;5��    M   .       	                	              �    M   /                                       �    M   .                                     �    M   .                                     �    M   .                                     5�_�                 N   3    ����                                                                                                                                                                                                                                                                                                                            =          =          v       f�   3 �   M   O   T      D            assert false report integer'image(HEXA*2) severity note;5��    M   3                                     �    M   4                                       �    M   3              	                	       �    M   3       	                	              �    M   3              	                	       5�_�                 >   5    ����                                                                                                                                                                                                                                                                                                                            =          =          v       f��     �   =   ?   U          �   =   ?   T    5��    =                      �                     �    =                  
   �              
       �    =                                          �    =                                        �    =                                          �    =                     
                     �    =                    	                    �    =                     
                     �    =                    	                    5�_�                 K       ����                                                                                                                                                                                                                                                                                                                            =          =          v       f��     �   K   M   V                  �   K   M   U    5��    K                                    	       �    K                                         �    K                     -                     �    K                     ,                     �    K                 	   +             	       �    K          	          +      	              �    K                 
   +             
       5�_�                   P   .    ����                                                                                                                                                                                                                                                                                                                            =          =          v       f�   4 �   O   Q   V      L            assert false report integer'image(HEXA*iteration) severity note;5��    O   .                 Q                    5�_�                 K       ����                                                                                                                                                                                                                                                                                                                            =          =          v       f��     �   J   L   R      S            w-- assert false report integer'image((iteration*16)+15) severity note;5��    J                     �                     5�_�  
                 
    ����                                                                                                                                                                                                                                                                                                                            =          =          v       f�_     �      !        5��                          �                     5�_�                   L   .    ����                                                                                                                                                                                                                                                                                                                            =          =          v       f�i   0 �   K   M   R      A            assert false report integer'image(2*3) severity note;5��    K   .                 �                    5�_�                 =       ����                                                                                                                                                                                                                                                                                                                            =          =   .       v       f��   / �   =   >   R    �   <   >   R      4    signal iteration: integer range -512 to 511:= 0;5��    <                    �                    5�_�  �  �         �   L        ����                                                                                                                                                                                                                                                                                                                            L   I       <           v        f�]     �   K   M   R      J            assert false report natural'image(iteration*16) severity note;5��    K                     �                    5�_�  �  �          �   8       ����                                                                                                                                                                                                                                                                                                                            L   I       <           v        f�h     �   7   9   R      F            count : out natural       -- 6-bit count output (64 steps)5��    7                    z                    5�_�  �  �          �   =       ����                                                                                                                                                                                                                                                                                                                            L   I       <           v        f�m     �   <   >   R      #    signal iteration: natural := 0;5��    <                    �                    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            L   I       <           v        f�z     �      	   R      B        count : out natural       -- 6-bit count output (64 steps)5��                        �                     5�_�  �              �          ����                                                                                                                                                                                                                                                                                                                            L   I       <           v        f��     �         R      !    count <= to_natural(counter);5��              
       
   l      
       
       5�_�  �  �      �  �   I   9    ����                                                                                                                                                                                                                                                                                                                            J   B       J   B       v   B    f�2   ' �   H   J   R      @            -- w <= msgi((iteration*16)+15 downto iteration*16);5��    H                     �      >       A       5�_�  �              �   J   9    ����                                                                                                                                                                                                                                                                                                                            J   B       J   B       v   B    f�A   ( �   I   K   R      X            -- assert false report integer'image(to_integer(unsigned(w))) severity note;5��    I                           V       Y       5�_�  �          �  �   I   #    ����                                                                                                                                                                                                                                                                                                                            J   B       J   B       v   B    f��     �   H   J   P      :            w <= msgi((iteration)+15 downto iteration*16);5��    H   "                  �                     �    H   !                  �                     �    H                      �                     5�_�  �  �      �  �   E       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��     �   D   F        5��    D                      �                     5�_�  �  �  �      �   F       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��     �   E   G        5��    E                      �                     5�_�  �              �   E       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��    �   D   F   I      Y        assert false report integer'image(to_integer(unsigned(iteration))) severity note;5��    D                     �                     5�_�  �          �  �   F       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��     �   E   G        5��    E                      �                     5�_�  �          �  �   <        ����                                                                                                                                                                                                                                                                                                                            #          &          V       f��     �   ;   >        5��    ;                      �      Z               5�_�  �  �      �  �   Q       ����                                                                                                                                                                                                                                                                                                                            T           O           V        fu     �   P   R        5��    P                            #               5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                            R          Q                 fu     �   R   T        5��    R                      �                     5�_�  �  �          �   Q       ����                                                                                                                                                                                                                                                                                                                            R          Q                 fu     �   P   R   V      "        wait for CLOCK_PERIOD / 2;5��    P                                          5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                            R          Q                 fu     �   Q   S   V      Y        assert false report integer'image(to_integer(unsigned(iteration))) severity note;5��    Q                     8                     5�_�  �  �          �   Q       ����                                                                                                                                                                                                                                                                                                                            R          Q                 fu     �   P   R   V              wait for CLOCK_PERIOD ;5��    P                     +                     5�_�  �  �          �   Q       ����                                                                                                                                                                                                                                                                                                                            R          Q                 fu     �   P   R   V              wait for CLOCK_PERIOD;5��    P                     *                     5�_�  �  �          �   Q       ����                                                                                                                                                                                                                                                                                                                            Q          Q                 fu     �   P   R        5��    P                                           5�_�  �  �          �   Q       ����                                                                                                                                                                                                                                                                                                                            Q          Q                 fu      �   Q   R   U    �   Q   R   U              wait for CLOCK_PERIOD;5��    Q                      g                     5�_�  �              �   R       ����                                                                                                                                                                                                                                                                                                                            Q          Q                 fu"    �   R   S   V    �   R   S   V      Y        assert false report integer'image(to_integer(unsigned(iteration))) severity note;5��    R                      �              Z       5�_�  �          �  �   q       ����                                                                                                                                                                                                                                                                                                                            �          q          V       fq    �   p   �   �          -- type h_vector is record   )    --     H_0 : bit_vector(31 downto 0);   )    --     H_1 : bit_vector(31 downto 0);   )    --     H_2 : bit_vector(31 downto 0);   )    --     H_3 : bit_vector(31 downto 0);   )    --     H_4 : bit_vector(31 downto 0);   )    --     H_5 : bit_vector(31 downto 0);   )    --     H_6 : bit_vector(31 downto 0);   )    --     H_7 : bit_vector(31 downto 0);       -- end record;       --   !    -- constant H : h_vector := (   <    --     H_0 => bit_vector(to_unsigned(32, 16#6a09e667#)),   <    --     H_1 => bit_vector(to_unsigned(32, 16#bb67ae85#)),   <    --     H_2 => bit_vector(to_unsigned(32, 16#3c6ef372#)),   <    --     H_3 => bit_vector(to_unsigned(32, 16#a54ff53a#)),   <    --     H_4 => bit_vector(to_unsigned(32, 16#510e527f#)),   <    --     H_5 => bit_vector(to_unsigned(32, 16#9b05688c#)),   <    --     H_6 => bit_vector(to_unsigned(32, 16#1f83d9ab#)),   ;    --     H_7 => bit_vector(to_unsigned(32, 16#5be0cd19#))   	    -- );5��    p                     �      Z      �      5�_�            �  �   /        ����                                                                                                                                                                                                                                                                                                                3           v          �   9          9    fp�     �   /   0   �    �   .   p   �   A   *bit_vector(to_unsigned(32, 16#428a2f98#)),   0bit_vector(to_unsigned(32, 16#71374491#)),    );   *bit_vector(to_unsigned(32, 16#b5c0fbcf#)),   Ebit_vector(to_unsigned(32, 16#e9b5dba5#)),    type k_vector is record   Pbit_vector(to_unsigned(32, 16#3956c25b#)),        K_0 : bit_vector(31 downto 0);   Pbit_vector(to_unsigned(32, 16#59f111f1#)),        K_1 : bit_vector(31 downto 0);   Pbit_vector(to_unsigned(32, 16#923f82a4#)),        K_2 : bit_vector(31 downto 0);   Pbit_vector(to_unsigned(32, 16#ab1c5ed5#)),        K_3 : bit_vector(31 downto 0);   Pbit_vector(to_unsigned(32, 16#d807aa98#)),        K_4 : bit_vector(31 downto 0);   Pbit_vector(to_unsigned(32, 16#12835b01#)),        K_5 : bit_vector(31 downto 0);   Pbit_vector(to_unsigned(32, 16#243185be#)),        K_6 : bit_vector(31 downto 0);   Pbit_vector(to_unsigned(32, 16#550c7dc3#)),        K_7 : bit_vector(31 downto 0);   Pbit_vector(to_unsigned(32, 16#72be5d74#)),        K_8 : bit_vector(31 downto 0);   Pbit_vector(to_unsigned(32, 16#80deb1fe#)),        K_9 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#9bdc06a7#)),        K_10 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#c19bf174#)),        K_11 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#e49b69c1#)),        K_12 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#efbe4786#)),        K_13 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#0fc19dc6#)),        K_14 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#240ca1cc#)),        K_15 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#2de92c6f#)),        K_16 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#4a7484aa#)),        K_17 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#5cb0a9dc#)),        K_18 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#76f988da#)),        K_19 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#983e5152#)),        K_20 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#a831c66d#)),        K_21 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#b00327c8#)),        K_22 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#bf597fc7#)),        K_23 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#c6e00bf3#)),        K_24 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#d5a79147#)),        K_25 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#06ca6351#)),        K_26 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#14292967#)),        K_27 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#27b70a85#)),        K_28 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#2e1b2138#)),        K_29 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#4d2c6dfc#)),        K_30 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#53380d13#)),        K_31 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#650a7354#)),        K_32 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#766a0abb#)),        K_33 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#81c2c92e#)),        K_34 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#92722c85#)),        K_35 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#a2bfe8a1#)),        K_36 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#a81a664b#)),        K_37 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#c24b8b70#)),        K_38 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#c76c51a3#)),        K_39 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#d192e819#)),        K_40 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#d6990624#)),        K_41 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#f40e3585#)),        K_42 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#106aa070#)),        K_43 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#19a4c116#)),        K_44 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#1e376c08#)),        K_45 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#2748774c#)),        K_46 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#34b0bcb5#)),        K_47 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#391c0cb3#)),        K_48 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#4ed8aa4a#)),        K_49 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#5b9cca4f#)),        K_50 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#682e6ff3#)),        K_51 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#748f82ee#)),        K_52 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#78a5636f#)),        K_53 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#84c87814#)),        K_54 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#8cc70208#)),        K_55 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#90befffa#)),        K_56 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#a4506ceb#)),        K_57 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#bef9a3f7#)),        K_58 : bit_vector(31 downto 0);   Qbit_vector(to_unsigned(32, 16#c67178f2#))         K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);5��    .                   *   )              *       �    /                   *   T              *       �    0                   *   �              *       �    1                   *   �              *       �    2                   *   �              *       �    3                   *   G              *       �    4                   *   �              *       �    5                   *   �              *       �    6                   *   :              *       �    7                   *   �              *       �    8                   *   �              *       �    9                   *   -              *       �    :                   *   ~              *       �    ;                   *   �              *       �    <                   *                  *       �    =                   *   r              *       �    >                   *   �              *       �    ?                   *   	              *       �    @                   *   h	              *       �    A                   *   �	              *       �    B                   *   
              *       �    C                   *   ^
              *       �    D                   *   �
              *       �    E                   *                 *       �    F                   *   T              *       �    G                   *   �              *       �    H                   *   �              *       �    I                   *   J              *       �    J                   *   �              *       �    K                   *   �              *       �    L                   *   @              *       �    M                   *   �              *       �    N                   *   �              *       �    O                   *   6              *       �    P                   *   �              *       �    Q                   *   �              *       �    R                   *   ,              *       �    S                   *   ~              *       �    T                   *   �              *       �    U                   *   "              *       �    V                   *   t              *       �    W                   *   �              *       �    X                   *                 *       �    Y                   *   j              *       �    Z                   *   �              *       �    [                   *                 *       �    \                   *   `              *       �    ]                   *   �              *       �    ^                   *                 *       �    _                   *   V              *       �    `                   *   �              *       �    a                   *   �              *       �    b                   *   L              *       �    c                   *   �              *       �    d                   *   �              *       �    e                   *   B              *       �    f                   *   �              *       �    g                   *   �              *       �    h                   *   8              *       �    i                   *   �              *       �    j                   *   �              *       �    k                   *   .              *       �    l                   *   �              *       �    m                   *   �              *       5�_�  }            ~   .       ����                                                                                                                                                                                                                                                                                                                2           u          �   9          9    fp�     �   .   /   �    �   -   o   �   A   F    signal k : k_bit_vector(to_unsigned(32, 16#428a2f98#)),vector := (   ;    );           bit_vector(to_unsigned(32, 16#71374491#)),   ;                 bit_vector(to_unsigned(32, 16#b5c0fbcf#)),   E    type k_vectorbit_vector(to_unsigned(32, 16#e9b5dba5#)), is record   P        K_0 : bitbit_vector(to_unsigned(32, 16#3956c25b#)),_vector(31 downto 0);   P        K_1 : bitbit_vector(to_unsigned(32, 16#59f111f1#)),_vector(31 downto 0);   P        K_2 : bitbit_vector(to_unsigned(32, 16#923f82a4#)),_vector(31 downto 0);   P        K_3 : bitbit_vector(to_unsigned(32, 16#ab1c5ed5#)),_vector(31 downto 0);   P        K_4 : bitbit_vector(to_unsigned(32, 16#d807aa98#)),_vector(31 downto 0);   P        K_5 : bitbit_vector(to_unsigned(32, 16#12835b01#)),_vector(31 downto 0);   P        K_6 : bitbit_vector(to_unsigned(32, 16#243185be#)),_vector(31 downto 0);   P        K_7 : bitbit_vector(to_unsigned(32, 16#550c7dc3#)),_vector(31 downto 0);   P        K_8 : bitbit_vector(to_unsigned(32, 16#72be5d74#)),_vector(31 downto 0);   P        K_9 : bitbit_vector(to_unsigned(32, 16#80deb1fe#)),_vector(31 downto 0);   Q        K_10 : bibit_vector(to_unsigned(32, 16#9bdc06a7#)),t_vector(31 downto 0);   Q        K_11 : bibit_vector(to_unsigned(32, 16#c19bf174#)),t_vector(31 downto 0);   Q        K_12 : bibit_vector(to_unsigned(32, 16#e49b69c1#)),t_vector(31 downto 0);   Q        K_13 : bibit_vector(to_unsigned(32, 16#efbe4786#)),t_vector(31 downto 0);   Q        K_14 : bibit_vector(to_unsigned(32, 16#0fc19dc6#)),t_vector(31 downto 0);   Q        K_15 : bibit_vector(to_unsigned(32, 16#240ca1cc#)),t_vector(31 downto 0);   Q        K_16 : bibit_vector(to_unsigned(32, 16#2de92c6f#)),t_vector(31 downto 0);   Q        K_17 : bibit_vector(to_unsigned(32, 16#4a7484aa#)),t_vector(31 downto 0);   Q        K_18 : bibit_vector(to_unsigned(32, 16#5cb0a9dc#)),t_vector(31 downto 0);   Q        K_19 : bibit_vector(to_unsigned(32, 16#76f988da#)),t_vector(31 downto 0);   Q        K_20 : bibit_vector(to_unsigned(32, 16#983e5152#)),t_vector(31 downto 0);   Q        K_21 : bibit_vector(to_unsigned(32, 16#a831c66d#)),t_vector(31 downto 0);   Q        K_22 : bibit_vector(to_unsigned(32, 16#b00327c8#)),t_vector(31 downto 0);   Q        K_23 : bibit_vector(to_unsigned(32, 16#bf597fc7#)),t_vector(31 downto 0);   Q        K_24 : bibit_vector(to_unsigned(32, 16#c6e00bf3#)),t_vector(31 downto 0);   Q        K_25 : bibit_vector(to_unsigned(32, 16#d5a79147#)),t_vector(31 downto 0);   Q        K_26 : bibit_vector(to_unsigned(32, 16#06ca6351#)),t_vector(31 downto 0);   Q        K_27 : bibit_vector(to_unsigned(32, 16#14292967#)),t_vector(31 downto 0);   Q        K_28 : bibit_vector(to_unsigned(32, 16#27b70a85#)),t_vector(31 downto 0);   Q        K_29 : bibit_vector(to_unsigned(32, 16#2e1b2138#)),t_vector(31 downto 0);   Q        K_30 : bibit_vector(to_unsigned(32, 16#4d2c6dfc#)),t_vector(31 downto 0);   Q        K_31 : bibit_vector(to_unsigned(32, 16#53380d13#)),t_vector(31 downto 0);   Q        K_32 : bibit_vector(to_unsigned(32, 16#650a7354#)),t_vector(31 downto 0);   Q        K_33 : bibit_vector(to_unsigned(32, 16#766a0abb#)),t_vector(31 downto 0);   Q        K_34 : bibit_vector(to_unsigned(32, 16#81c2c92e#)),t_vector(31 downto 0);   Q        K_35 : bibit_vector(to_unsigned(32, 16#92722c85#)),t_vector(31 downto 0);   Q        K_36 : bibit_vector(to_unsigned(32, 16#a2bfe8a1#)),t_vector(31 downto 0);   Q        K_37 : bibit_vector(to_unsigned(32, 16#a81a664b#)),t_vector(31 downto 0);   Q        K_38 : bibit_vector(to_unsigned(32, 16#c24b8b70#)),t_vector(31 downto 0);   Q        K_39 : bibit_vector(to_unsigned(32, 16#c76c51a3#)),t_vector(31 downto 0);   Q        K_40 : bibit_vector(to_unsigned(32, 16#d192e819#)),t_vector(31 downto 0);   Q        K_41 : bibit_vector(to_unsigned(32, 16#d6990624#)),t_vector(31 downto 0);   Q        K_42 : bibit_vector(to_unsigned(32, 16#f40e3585#)),t_vector(31 downto 0);   Q        K_43 : bibit_vector(to_unsigned(32, 16#106aa070#)),t_vector(31 downto 0);   Q        K_44 : bibit_vector(to_unsigned(32, 16#19a4c116#)),t_vector(31 downto 0);   Q        K_45 : bibit_vector(to_unsigned(32, 16#1e376c08#)),t_vector(31 downto 0);   Q        K_46 : bibit_vector(to_unsigned(32, 16#2748774c#)),t_vector(31 downto 0);   Q        K_47 : bibit_vector(to_unsigned(32, 16#34b0bcb5#)),t_vector(31 downto 0);   Q        K_48 : bibit_vector(to_unsigned(32, 16#391c0cb3#)),t_vector(31 downto 0);   Q        K_49 : bibit_vector(to_unsigned(32, 16#4ed8aa4a#)),t_vector(31 downto 0);   Q        K_50 : bibit_vector(to_unsigned(32, 16#5b9cca4f#)),t_vector(31 downto 0);   Q        K_51 : bibit_vector(to_unsigned(32, 16#682e6ff3#)),t_vector(31 downto 0);   Q        K_52 : bibit_vector(to_unsigned(32, 16#748f82ee#)),t_vector(31 downto 0);   Q        K_53 : bibit_vector(to_unsigned(32, 16#78a5636f#)),t_vector(31 downto 0);   Q        K_54 : bibit_vector(to_unsigned(32, 16#84c87814#)),t_vector(31 downto 0);   Q        K_55 : bibit_vector(to_unsigned(32, 16#8cc70208#)),t_vector(31 downto 0);   Q        K_56 : bibit_vector(to_unsigned(32, 16#90befffa#)),t_vector(31 downto 0);   Q        K_57 : bibit_vector(to_unsigned(32, 16#a4506ceb#)),t_vector(31 downto 0);   Q        K_58 : bibit_vector(to_unsigned(32, 16#bef9a3f7#)),t_vector(31 downto 0);   Q        K_59 : bibit_vector(to_unsigned(32, 16#c67178f2#)) t_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);5��    -                  *                 *       �    .                  5   Y              5       �    /                   ;   �              ;       �    0                  *   �              *       �    1                  *   "              *       �    2                  *   s              *       �    3                  *   �              *       �    4                  *                 *       �    5                  *   f              *       �    6                  *   �              *       �    7                  *                 *       �    8                  *   Y              *       �    9                  *   �              *       �    :                  *   �              *       �    ;                  *   L              *       �    <                  *   �              *       �    =                  *   �              *       �    >                  *   B	              *       �    ?                  *   �	              *       �    @                  *   �	              *       �    A                  *   8
              *       �    B                  *   �
              *       �    C                  *   �
              *       �    D                  *   .              *       �    E                  *   �              *       �    F                  *   �              *       �    G                  *   $              *       �    H                  *   v              *       �    I                  *   �              *       �    J                  *                 *       �    K                  *   l              *       �    L                  *   �              *       �    M                  *                 *       �    N                  *   b              *       �    O                  *   �              *       �    P                  *                 *       �    Q                  *   X              *       �    R                  *   �              *       �    S                  *   �              *       �    T                  *   N              *       �    U                  *   �              *       �    V                  *   �              *       �    W                  *   D              *       �    X                  *   �              *       �    Y                  *   �              *       �    Z                  *   :              *       �    [                  *   �              *       �    \                  *   �              *       �    ]                  *   0              *       �    ^                  *   �              *       �    _                  *   �              *       �    `                  *   &              *       �    a                  *   x              *       �    b                  *   �              *       �    c                  *                 *       �    d                  *   n              *       �    e                  *   �              *       �    f                  *                 *       �    g                  *   d              *       �    h                  *   �              *       �    i                  *                 *       �    j                  *   Z              *       �    k                  *   �              *       �    l                  *   �              *       5�_�  z          |  {   /       ����                                                                                                                                                                                                                                                                                                                6           /          n   -          -    fp�     �   .   3   �                                  �   /   0   �    �   .   p   �   A   /    bit_vector(to_unsigned(32, 16#428a2f98#)),    /    bit_vector(to_unsigned(32, 16#71374491#)),    /    bit_vector(to_unsigned(32, 16#b5c0fbcf#)),    .    bit_vector(to_unsigned(32, 16#e9b5dba5#)),   0    bit_vector(to_unsigned(32, 16#3956c25b#)),);   .    bit_vector(to_unsigned(32, 16#59f111f1#)),   E    bit_vector(to_unsigned(32, 16#923f82a4#)),type k_vector is record   P    bit_vector(to_unsigned(32, 16#ab1c5ed5#)),    K_0 : bit_vector(31 downto 0);   P    bit_vector(to_unsigned(32, 16#d807aa98#)),    K_1 : bit_vector(31 downto 0);   P    bit_vector(to_unsigned(32, 16#12835b01#)),    K_2 : bit_vector(31 downto 0);   P    bit_vector(to_unsigned(32, 16#243185be#)),    K_3 : bit_vector(31 downto 0);   P    bit_vector(to_unsigned(32, 16#550c7dc3#)),    K_4 : bit_vector(31 downto 0);   P    bit_vector(to_unsigned(32, 16#72be5d74#)),    K_5 : bit_vector(31 downto 0);   P    bit_vector(to_unsigned(32, 16#80deb1fe#)),    K_6 : bit_vector(31 downto 0);   P    bit_vector(to_unsigned(32, 16#9bdc06a7#)),    K_7 : bit_vector(31 downto 0);   P    bit_vector(to_unsigned(32, 16#c19bf174#)),    K_8 : bit_vector(31 downto 0);   P    bit_vector(to_unsigned(32, 16#e49b69c1#)),    K_9 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#efbe4786#)),    K_10 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#0fc19dc6#)),    K_11 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#240ca1cc#)),    K_12 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#2de92c6f#)),    K_13 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#4a7484aa#)),    K_14 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#5cb0a9dc#)),    K_15 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#76f988da#)),    K_16 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#983e5152#)),    K_17 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#a831c66d#)),    K_18 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#b00327c8#)),    K_19 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#bf597fc7#)),    K_20 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#c6e00bf3#)),    K_21 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#d5a79147#)),    K_22 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#06ca6351#)),    K_23 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#14292967#)),    K_24 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#27b70a85#)),    K_25 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#2e1b2138#)),    K_26 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#4d2c6dfc#)),    K_27 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#53380d13#)),    K_28 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#650a7354#)),    K_29 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#766a0abb#)),    K_30 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#81c2c92e#)),    K_31 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#92722c85#)),    K_32 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#a2bfe8a1#)),    K_33 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#a81a664b#)),    K_34 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#c24b8b70#)),    K_35 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#c76c51a3#)),    K_36 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#d192e819#)),    K_37 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#d6990624#)),    K_38 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#f40e3585#)),    K_39 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#106aa070#)),    K_40 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#19a4c116#)),    K_41 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#1e376c08#)),    K_42 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#2748774c#)),    K_43 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#34b0bcb5#)),    K_44 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#391c0cb3#)),    K_45 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#4ed8aa4a#)),    K_46 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#5b9cca4f#)),    K_47 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#682e6ff3#)),    K_48 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#748f82ee#)),    K_49 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#78a5636f#)),    K_50 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#84c87814#)),    K_51 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#8cc70208#)),    K_52 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#90befffa#)),    K_53 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#a4506ceb#)),    K_54 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#bef9a3f7#)),    K_55 : bit_vector(31 downto 0);   Q    bit_vector(to_unsigned(32, 16#c67178f2#))     K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);5��    .          *           -      *               �    /          *           3      *               �    0          *           9      *               �    1          )           ?      )               �    .                  *   -              *       �    /                  *   ]              *       �    0                  *   �              *       �    1                  *   �              *       �    2                  *   �              *       �    3                   .                 .       �    4                  *   L              *       �    5                  *   �              *       �    6                  *   �              *       �    7                  *   4              *       �    8                  *   �              *       �    9                  *   �              *       �    :                  *   '              *       �    ;                  *   x              *       �    <                  *   �              *       �    =                  *                 *       �    >                  *   k              *       �    ?                  *   �              *       �    @                  *   	              *       �    A                  *   `	              *       �    B                  *   �	              *       �    C                  *   
              *       �    D                  *   V
              *       �    E                  *   �
              *       �    F                  *   �
              *       �    G                  *   L              *       �    H                  *   �              *       �    I                  *   �              *       �    J                  *   B              *       �    K                  *   �              *       �    L                  *   �              *       �    M                  *   8              *       �    N                  *   �              *       �    O                  *   �              *       �    P                  *   .              *       �    Q                  *   �              *       �    R                  *   �              *       �    S                  *   $              *       �    T                  *   v              *       �    U                  *   �              *       �    V                  *                 *       �    W                  *   l              *       �    X                  *   �              *       �    Y                  *                 *       �    Z                  *   b              *       �    [                  *   �              *       �    \                  *                 *       �    ]                  *   X              *       �    ^                  *   �              *       �    _                  *   �              *       �    `                  *   N              *       �    a                  *   �              *       �    b                  *   �              *       �    c                  *   D              *       �    d                  *   �              *       �    e                  *   �              *       �    f                  *   :              *       �    g                  *   �              *       �    h                  *   �              *       �    i                  *   0              *       �    j                  *   �              *       �    k                  *   �              *       �    l                  *   &              *       �    m                  *   x              *       5�_�  m          o  n   -   '    ����                                                                                                                                                                                                                                                                                                                1           .          .          v       fp     �   ,   .   �      (    type k_vector is array(0 to 63) of ;5��    ,   '                  �                     5�_�  e          g  f          ����                                                                                                                                                                                                                                                                                                                -           p          �          V       fnz     �               5��                          �                     5�_�  O          Q  P           ����                                                                                                                                                                                                                                                                                                                            �          �           V       fP     �              5��                                                5�_�  ,  .      M  -   >       ����                                                                                                                                                                                                                                                                                                                >           �          =          V       f�     �   <   =   �   �       -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );              type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   7        H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   7        H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   7        H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   7        H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   7        H_4 => bit_vector(to_signed(32, 16#510e527f#)),   7        H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   7        H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   6        H_7 => bit_vector(to_signed(32, 16#5be0cd19#))       );�   �  v      �   <   �       �       -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))       );5��   =       �       <       )      �      (      �    �                     {                    �    �                     �                    �    �                     �                    �    �                                         �    �                     K                    �    �                                         �    �                     �                    �    �                     �                    �    �                                         �    �                     O                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     "                    �    �                     W                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     +                    �    �                     `                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     4                    �    �                     i                    �    �                     �                    �    �                     �                    �    �                                         �    �                     =                    �    �                     r                    �    �                     �                    �    �                     �                    �    �                                         �    �                     F                    �    �                     {                    �    �                     �                    �    �                     �                    �    �                                         �    �                     O                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     #                    �    �                     X                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     ,                    �    �                     a                    �    �                     �                    �    �                     �                    �    �                                          �    �                     5                    �    �                     j                    �    �                     �                    �    �                     �                    �    �                     	                    �    �                     >                    �    �                     s                    �    �                     �                    �    �                     �                    �    �                                         �    �                     G                    �    �                     |                    �    �                      �                     �    �                      �                     �    �                      �                     �    �                     �                    �    �                     �                    �    �                                         �    �                     5                    �    �                     X                    �    �                     {                    �    �                     �                    �    �                     �                    �    �                      �                     �    �                      �                     �    �                                           �    �                      <                     �    �                      l                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      ,                      �    �                      \                      5�_�  -  /          .   =       ����                                                                                                                                                                                                                                                                                                                =           �          <          V       f�     �   ;   <   �   �       -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))       );�   �  u      �   ;   �       �       -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   <       �       ;       (      j            �    <                     &                    �    =                     F                    �    >                     q                    �    ?                     �                    �    @                     �                    �    A                     �                    �    B                                         �    C                     H                    �    D                     s                    �    E                     �                    �    F                     �                    �    G                     �                    �    H                                          �    I                     L                    �    J                     x                    �    K                     �                    �    L                     �                    �    M                     �                    �    N                     (	                    �    O                     T	                    �    P                     �	                    �    Q                     �	                    �    R                     �	                    �    S                     
                    �    T                     0
                    �    U                     \
                    �    V                     �
                    �    W                     �
                    �    X                     �
                    �    Y                                         �    Z                     8                    �    [                     d                    �    \                     �                    �    ]                     �                    �    ^                     �                    �    _                                         �    `                     @                    �    a                     l                    �    b                     �                    �    c                     �                    �    d                     �                    �    e                                         �    f                     H                    �    g                     t                    �    h                     �                    �    i                     �                    �    j                     �                    �    k                     $                    �    l                     P                    �    m                     |                    �    n                     �                    �    o                     �                    �    p                                          �    q                     ,                    �    r                     X                    �    s                     �                    �    t                     �                    �    u                     �                    �    v                                         �    w                     4                    �    x                     `                    �    y                     �                    �    z                     �                    �    {                     �                    �    |                                         �    }                     <                    �                         Q                    �    �                     t                    �    �                     �                    �    �                     �                    �    �                                         �    �                     T                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     4                    �    �                     l                    �    �                     �                    �    �                     �                    �    �                                         �    �                     O                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     3                    �    �                     l                    �    �                     �                    �    �                     �                    �    �                                         �    �                     P                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     4                    �    �                     m                    �    �                     �                    �    �                     �                    �    �                                         �    �                     Q                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     5                    �    �                     n                    �    �                     �                    �    �                     �                    �    �                                         �    �                     R                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     6                    �    �                     o                    �    �                     �                    �    �                     �                    �    �                                         �    �                     S                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     7                    �    �                     p                    �    �                     �                    �    �                     �                    �    �                                         �    �                     T                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     8                    �    �                     q                    �    �                      �                     �    �                      �                     �    �                     �                    �    �                     �                    �    �                                          �    �                     B                     �    �                     i                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                      !                     �    �                      !                     �    �                      5!                     �    �                      i!                     �    �                      �!                     �    �                      �!                     �    �                      "                     �    �                      9"                     �    �                      m"                     �    �                      �"                     �    �                      �"                     5�_�  .  0          /   <       ����                                                                                                                                                                                                                                                                                                                <           �          ;          V       f�     �   :   ;   �   �       -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  t      �   :   �       �   A                                                     -- Constants   #            type k_vector is record   .                K_0 : bit_vector(31 downto 0);   .                K_1 : bit_vector(31 downto 0);   .                K_2 : bit_vector(31 downto 0);   .                K_3 : bit_vector(31 downto 0);   .                K_4 : bit_vector(31 downto 0);   .                K_5 : bit_vector(31 downto 0);   .                K_6 : bit_vector(31 downto 0);   .                K_7 : bit_vector(31 downto 0);   .                K_8 : bit_vector(31 downto 0);   .                K_9 : bit_vector(31 downto 0);   /                K_10 : bit_vector(31 downto 0);   /                K_11 : bit_vector(31 downto 0);   /                K_12 : bit_vector(31 downto 0);   /                K_13 : bit_vector(31 downto 0);   /                K_14 : bit_vector(31 downto 0);   /                K_15 : bit_vector(31 downto 0);   /                K_16 : bit_vector(31 downto 0);   /                K_17 : bit_vector(31 downto 0);   /                K_18 : bit_vector(31 downto 0);   /                K_19 : bit_vector(31 downto 0);   /                K_20 : bit_vector(31 downto 0);   /                K_21 : bit_vector(31 downto 0);   /                K_22 : bit_vector(31 downto 0);   /                K_23 : bit_vector(31 downto 0);   /                K_24 : bit_vector(31 downto 0);   /                K_25 : bit_vector(31 downto 0);   /                K_26 : bit_vector(31 downto 0);   /                K_27 : bit_vector(31 downto 0);   /                K_28 : bit_vector(31 downto 0);   /                K_29 : bit_vector(31 downto 0);   /                K_30 : bit_vector(31 downto 0);   /                K_31 : bit_vector(31 downto 0);   /                K_32 : bit_vector(31 downto 0);   /                K_33 : bit_vector(31 downto 0);   /                K_34 : bit_vector(31 downto 0);   /                K_35 : bit_vector(31 downto 0);   /                K_36 : bit_vector(31 downto 0);   /                K_37 : bit_vector(31 downto 0);   /                K_38 : bit_vector(31 downto 0);   /                K_39 : bit_vector(31 downto 0);   /                K_40 : bit_vector(31 downto 0);   /                K_41 : bit_vector(31 downto 0);   /                K_42 : bit_vector(31 downto 0);   /                K_43 : bit_vector(31 downto 0);   /                K_44 : bit_vector(31 downto 0);   /                K_45 : bit_vector(31 downto 0);   /                K_46 : bit_vector(31 downto 0);   /                K_47 : bit_vector(31 downto 0);   /                K_48 : bit_vector(31 downto 0);   /                K_49 : bit_vector(31 downto 0);   /                K_50 : bit_vector(31 downto 0);   /                K_51 : bit_vector(31 downto 0);   /                K_52 : bit_vector(31 downto 0);   /                K_53 : bit_vector(31 downto 0);   /                K_54 : bit_vector(31 downto 0);   /                K_55 : bit_vector(31 downto 0);   /                K_56 : bit_vector(31 downto 0);   /                K_57 : bit_vector(31 downto 0);   /                K_58 : bit_vector(31 downto 0);   /                K_59 : bit_vector(31 downto 0);   /                K_60 : bit_vector(31 downto 0);   /                K_61 : bit_vector(31 downto 0);   /                K_62 : bit_vector(31 downto 0);   /                K_63 : bit_vector(31 downto 0);               end record;       &            constant K : k_vector := (   ;            K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   ;            K_1 => bit_vector(to_signed(32, 16#71374491#)),   ;            K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   ;            K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   ;            K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   ;            K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   ;            K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   ;            K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   ;            K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   ;            K_9 => bit_vector(to_signed(32, 16#12835b01#)),   <            K_10 => bit_vector(to_signed(32, 16#243185be#)),   <            K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   <            K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   <            K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   <            K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   <            K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   <            K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   <            K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   <            K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   <            K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   <            K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   <            K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   <            K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   <            K_23 => bit_vector(to_signed(32, 16#76f988da#)),   <            K_24 => bit_vector(to_signed(32, 16#983e5152#)),   <            K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   <            K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   <            K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   <            K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   <            K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   <            K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   <            K_31 => bit_vector(to_signed(32, 16#14292967#)),   <            K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   <            K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   <            K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   <            K_35 => bit_vector(to_signed(32, 16#53380d13#)),   <            K_36 => bit_vector(to_signed(32, 16#650a7354#)),   <            K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   <            K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   <            K_39 => bit_vector(to_signed(32, 16#92722c85#)),   <            K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   <            K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   <            K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   <            K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   <            K_44 => bit_vector(to_signed(32, 16#d192e819#)),   <            K_45 => bit_vector(to_signed(32, 16#d6990624#)),   <            K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   <            K_47 => bit_vector(to_signed(32, 16#106aa070#)),   <            K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   <            K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   <            K_50 => bit_vector(to_signed(32, 16#2748774c#)),   <            K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   <            K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   <            K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   <            K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   <            K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   <            K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   <            K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   <            K_58 => bit_vector(to_signed(32, 16#84c87814#)),   <            K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   <            K_60 => bit_vector(to_signed(32, 16#90befffa#)),   <            K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   <            K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   ;            K_63 => bit_vector(to_signed(32, 16#c67178f2#))   
        );               type h_vector is record   *            H_0 : bit_vector(31 downto 0);   *            H_1 : bit_vector(31 downto 0);   *            H_2 : bit_vector(31 downto 0);   *            H_3 : bit_vector(31 downto 0);   *            H_4 : bit_vector(31 downto 0);   *            H_5 : bit_vector(31 downto 0);   *            H_6 : bit_vector(31 downto 0);   *            H_7 : bit_vector(31 downto 0);           end record;       "        constant H : h_vector := (   7        H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   7        H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   7        H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   7        H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   7        H_4 => bit_vector(to_signed(32, 16#510e527f#)),   7        H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   7        H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   6        H_7 => bit_vector(to_signed(32, 16#5be0cd19#))       );5��   ;       �       :             �      
      �    :                  5   
             5       �    ;                     L                    �    <                     p                    �    =                     �                    �    >                     �                    �    ?                     �                    �    @                     ,                    �    A                     [                    �    B                     �                    �    C                     �                    �    D                     �                    �    E                                         �    F                     F                    �    G                     v                    �    H                     �                    �    I                     �                    �    J                     	                    �    K                     6	                    �    L                     f	                    �    M                     �	                    �    N                     �	                    �    O                     �	                    �    P                     &
                    �    Q                     V
                    �    R                     �
                    �    S                     �
                    �    T                     �
                    �    U                                         �    V                     F                    �    W                     v                    �    X                     �                    �    Y                     �                    �    Z                                         �    [                     6                    �    \                     f                    �    ]                     �                    �    ^                     �                    �    _                     �                    �    `                     &                    �    a                     V                    �    b                     �                    �    c                     �                    �    d                     �                    �    e                                         �    f                     F                    �    g                     v                    �    h                     �                    �    i                     �                    �    j                                         �    k                     6                    �    l                     f                    �    m                     �                    �    n                     �                    �    o                     �                    �    p                     &                    �    q                     V                    �    r                     �                    �    s                     �                    �    t                     �                    �    u                                         �    v                     F                    �    w                     v                    �    x                     �                    �    y                     �                    �    z                                         �    {                     6                    �    |                     f                    �    ~                                         �                         �                    �    �                     �                    �    �                                         �    �                     Z                    �    �                     �                    �    �                     �                    �    �                                         �    �                     J                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     ;                    �    �                     x                    �    �                     �                    �    �                     �                    �    �                     /                    �    �                     l                    �    �                     �                    �    �                     �                    �    �                     #                    �    �                     `                    �    �                     �                    �    �                     �                    �    �                                         �    �                     T                    �    �                     �                    �    �                     �                    �    �                                         �    �                     H                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     <                    �    �                     y                    �    �                     �                    �    �                     �                    �    �                     0                    �    �                     m                    �    �                     �                    �    �                     �                    �    �                     $                    �    �                     a                    �    �                     �                    �    �                     �                    �    �                                         �    �                     U                    �    �                     �                    �    �                     �                    �    �                                         �    �                     I                    �    �                     �                    �    �                     �                    �    �                                          �    �                     =                    �    �                     z                    �    �                     �                    �    �                     �                    �    �                     1                     �    �                     n                     �    �                     �                     �    �                     �                     �    �                     %!                    �    �                     b!                    �    �                     �!                    �    �                     �!                    �    �                     �!                    �    �                     "                    �    �                     2"                    �    �                     ]"                    �    �                     �"                    �    �                     �"                    �    �                     �"                    �    �                     	#                    �    �                     4#                    �    �                     _#                    �    �                     t#                    �    �                     �#                    �    �                     �#                    �    �                     $                    �    �                     ?$                    �    �                     w$                    �    �                     �$                    �    �                     �$                    �    �                     %                    �    �                      V%                     5�_�  /  1          0   ;       ����                                                                                                                                                                                                                                                                                                                ;           �          :          V       f�     �   9   :   �   �   A                                                     -- Constants   #            type k_vector is record   .                K_0 : bit_vector(31 downto 0);   .                K_1 : bit_vector(31 downto 0);   .                K_2 : bit_vector(31 downto 0);   .                K_3 : bit_vector(31 downto 0);   .                K_4 : bit_vector(31 downto 0);   .                K_5 : bit_vector(31 downto 0);   .                K_6 : bit_vector(31 downto 0);   .                K_7 : bit_vector(31 downto 0);   .                K_8 : bit_vector(31 downto 0);   .                K_9 : bit_vector(31 downto 0);   /                K_10 : bit_vector(31 downto 0);   /                K_11 : bit_vector(31 downto 0);   /                K_12 : bit_vector(31 downto 0);   /                K_13 : bit_vector(31 downto 0);   /                K_14 : bit_vector(31 downto 0);   /                K_15 : bit_vector(31 downto 0);   /                K_16 : bit_vector(31 downto 0);   /                K_17 : bit_vector(31 downto 0);   /                K_18 : bit_vector(31 downto 0);   /                K_19 : bit_vector(31 downto 0);   /                K_20 : bit_vector(31 downto 0);   /                K_21 : bit_vector(31 downto 0);   /                K_22 : bit_vector(31 downto 0);   /                K_23 : bit_vector(31 downto 0);   /                K_24 : bit_vector(31 downto 0);   /                K_25 : bit_vector(31 downto 0);   /                K_26 : bit_vector(31 downto 0);   /                K_27 : bit_vector(31 downto 0);   /                K_28 : bit_vector(31 downto 0);   /                K_29 : bit_vector(31 downto 0);   /                K_30 : bit_vector(31 downto 0);   /                K_31 : bit_vector(31 downto 0);   /                K_32 : bit_vector(31 downto 0);   /                K_33 : bit_vector(31 downto 0);   /                K_34 : bit_vector(31 downto 0);   /                K_35 : bit_vector(31 downto 0);   /                K_36 : bit_vector(31 downto 0);   /                K_37 : bit_vector(31 downto 0);   /                K_38 : bit_vector(31 downto 0);   /                K_39 : bit_vector(31 downto 0);   /                K_40 : bit_vector(31 downto 0);   /                K_41 : bit_vector(31 downto 0);   /                K_42 : bit_vector(31 downto 0);   /                K_43 : bit_vector(31 downto 0);   /                K_44 : bit_vector(31 downto 0);   /                K_45 : bit_vector(31 downto 0);   /                K_46 : bit_vector(31 downto 0);   /                K_47 : bit_vector(31 downto 0);   /                K_48 : bit_vector(31 downto 0);   /                K_49 : bit_vector(31 downto 0);   /                K_50 : bit_vector(31 downto 0);   /                K_51 : bit_vector(31 downto 0);   /                K_52 : bit_vector(31 downto 0);   /                K_53 : bit_vector(31 downto 0);   /                K_54 : bit_vector(31 downto 0);   /                K_55 : bit_vector(31 downto 0);   /                K_56 : bit_vector(31 downto 0);   /                K_57 : bit_vector(31 downto 0);   /                K_58 : bit_vector(31 downto 0);   /                K_59 : bit_vector(31 downto 0);   /                K_60 : bit_vector(31 downto 0);   /                K_61 : bit_vector(31 downto 0);   /                K_62 : bit_vector(31 downto 0);   /                K_63 : bit_vector(31 downto 0);               end record;       &            constant K : k_vector := (   ;            K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   ;            K_1 => bit_vector(to_signed(32, 16#71374491#)),   ;            K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   ;            K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   ;            K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   ;            K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   ;            K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   ;            K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   ;            K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   ;            K_9 => bit_vector(to_signed(32, 16#12835b01#)),   <            K_10 => bit_vector(to_signed(32, 16#243185be#)),   <            K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   <            K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   <            K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   <            K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   <            K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   <            K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   <            K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   <            K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   <            K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   <            K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   <            K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   <            K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   <            K_23 => bit_vector(to_signed(32, 16#76f988da#)),   <            K_24 => bit_vector(to_signed(32, 16#983e5152#)),   <            K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   <            K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   <            K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   <            K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   <            K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   <            K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   <            K_31 => bit_vector(to_signed(32, 16#14292967#)),   <            K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   <            K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   <            K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   <            K_35 => bit_vector(to_signed(32, 16#53380d13#)),   <            K_36 => bit_vector(to_signed(32, 16#650a7354#)),   <            K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   <            K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   <            K_39 => bit_vector(to_signed(32, 16#92722c85#)),   <            K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   <            K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   <            K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   <            K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   <            K_44 => bit_vector(to_signed(32, 16#d192e819#)),   <            K_45 => bit_vector(to_signed(32, 16#d6990624#)),   <            K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   <            K_47 => bit_vector(to_signed(32, 16#106aa070#)),   <            K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   <            K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   <            K_50 => bit_vector(to_signed(32, 16#2748774c#)),   <            K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   <            K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   <            K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   <            K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   <            K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   <            K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   <            K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   <            K_58 => bit_vector(to_signed(32, 16#84c87814#)),   <            K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   <            K_60 => bit_vector(to_signed(32, 16#90befffa#)),   <            K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   <            K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   ;            K_63 => bit_vector(to_signed(32, 16#c67178f2#))   
        );               type h_vector is record   *            H_0 : bit_vector(31 downto 0);   *            H_1 : bit_vector(31 downto 0);   *            H_2 : bit_vector(31 downto 0);   *            H_3 : bit_vector(31 downto 0);   *            H_4 : bit_vector(31 downto 0);   *            H_5 : bit_vector(31 downto 0);   *            H_6 : bit_vector(31 downto 0);   *            H_7 : bit_vector(31 downto 0);           end record;       "        constant H : h_vector := (   7        H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   7        H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   7        H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   7        H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   7        H_4 => bit_vector(to_signed(32, 16#510e527f#)),   7        H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   7        H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   6        H_7 => bit_vector(to_signed(32, 16#5be0cd19#))       );�   �  s      �   9   �       �   ?                                                   -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   :       �       9       
      S      �      �    9           5       3   �      5       3       �    :                     �                    �    ;                                         �    <                     ?                    �    =                     j                    �    >                     �                    �    ?                     �                    �    @                     �                    �    A                                         �    B                     A                    �    C                     l                    �    D                     �                    �    E                     �                    �    F                     �                    �    G                                         �    H                     F                    �    I                     r                    �    J                     �                    �    K                     �                    �    L                     �                    �    M                     "	                    �    N                     N	                    �    O                     z	                    �    P                     �	                    �    Q                     �	                    �    R                     �	                    �    S                     *
                    �    T                     V
                    �    U                     �
                    �    V                     �
                    �    W                     �
                    �    X                                         �    Y                     2                    �    Z                     ^                    �    [                     �                    �    \                     �                    �    ]                     �                    �    ^                                         �    _                     :                    �    `                     f                    �    a                     �                    �    b                     �                    �    c                     �                    �    d                                         �    e                     B                    �    f                     n                    �    g                     �                    �    h                     �                    �    i                     �                    �    j                                         �    k                     J                    �    l                     v                    �    m                     �                    �    n                     �                    �    o                     �                    �    p                     &                    �    q                     R                    �    r                     ~                    �    s                     �                    �    t                     �                    �    u                                         �    v                     .                    �    w                     Z                    �    x                     �                    �    y                     �                    �    z                     �                    �    {                     
                    �    }                                         �    ~                     B                    �                         z                    �    �                     �                    �    �                     �                    �    �                     "                    �    �                     Z                    �    �                     �                    �    �                     �                    �    �                                         �    �                     :                    �    �                     r                    �    �                     �                    �    �                     �                    �    �                                         �    �                     V                    �    �                     �                    �    �                     �                    �    �                                         �    �                     :                    �    �                     s                    �    �                     �                    �    �                     �                    �    �                                         �    �                     W                    �    �                     �                    �    �                     �                    �    �                                         �    �                     ;                    �    �                     t                    �    �                     �                    �    �                     �                    �    �                                         �    �                     X                    �    �                     �                    �    �                     �                    �    �                                         �    �                     <                    �    �                     u                    �    �                     �                    �    �                     �                    �    �                                          �    �                     Y                    �    �                     �                    �    �                     �                    �    �                                         �    �                     =                    �    �                     v                    �    �                     �                    �    �                     �                    �    �                     !                    �    �                     Z                    �    �                     �                    �    �                     �                    �    �                                         �    �                     >                    �    �                     w                    �    �                     �                    �    �                     �                    �    �                     "                    �    �                     [                    �    �                     �                    �    �                     �                    �    �                                         �    �                     ?                    �    �                     w                    �    �                                         �    �                     �                    �    �                     �                    �    �                     �                    �    �                                          �    �                     7                     �    �                     ^                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     !                    �    �                     7!                    �    �                     k!                    �    �                     �!                    �    �                     �!                    �    �                     "                    �    �                     ;"                    �    �                     o"                    �    �                      �"                     5�_�  0  2          1   :       ����                                                                                                                                                                                                                                                                                                                :           �          9          V       f�     �   8   9   �   �   ?                                                   -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  r      �   8   �       �   A                                                     -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   9       �       8       �      �      r      �    8           3       5   r      3       5       5�_�  1  3          2   9       ����                                                                                                                                                                                                                                                                                                                9           �          8          V       f�     �   7   8   �   �   A                                                     -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  q      �   7   �       �           -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   8       �       7       r      �      .      �    7           5          .      5              5�_�  2  4          3   8       ����                                                                                                                                                                                                                                                                                                                8           �          7          V       f�     �   6   7   �   �           -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  p      �   6   �       �           -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   7       �       6       .      �            �    7                     4                    �    8                     P                    �    9                     w                    �    :                     �                    �    ;                     �                    �    <                     �                    �    =                                         �    >                     :                    �    ?                     a                    �    @                     �                    �    A                     �                    �    B                     �                    �    C                     �                    �    D                     &                    �    E                     N                    �    F                     v                    �    G                     �                    �    H                     �                    �    I                     �                    �    J                                         �    K                     >                    �    L                     f                    �    M                     �                    �    N                     �                    �    O                     �                    �    P                     	                    �    Q                     .	                    �    R                     V	                    �    S                     ~	                    �    T                     �	                    �    U                     �	                    �    V                     �	                    �    W                     
                    �    X                     F
                    �    Y                     n
                    �    Z                     �
                    �    [                     �
                    �    \                     �
                    �    ]                                         �    ^                     6                    �    _                     ^                    �    `                     �                    �    a                     �                    �    b                     �                    �    c                     �                    �    d                     &                    �    e                     N                    �    f                     v                    �    g                     �                    �    h                     �                    �    i                     �                    �    j                                         �    k                     >                    �    l                     f                    �    m                     �                    �    n                     �                    �    o                     �                    �    p                                         �    q                     .                    �    r                     V                    �    s                     ~                    �    t                     �                    �    u                     �                    �    v                     �                    �    w                                         �    x                     F                    �    z                     W                    �    {                     v                    �    |                     �                    �    }                     �                    �    ~                                         �                         F                    �    �                     z                    �    �                     �                    �    �                     �                    �    �                                         �    �                     J                    �    �                     ~                    �    �                     �                    �    �                     �                    �    �                                         �    �                     R                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     &                    �    �                     [                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     /                    �    �                     d                    �    �                     �                    �    �                     �                    �    �                                         �    �                     8                    �    �                     m                    �    �                     �                    �    �                     �                    �    �                                         �    �                     A                    �    �                     v                    �    �                     �                    �    �                     �                    �    �                                         �    �                     J                    �    �                                         �    �                     �                    �    �                     �                    �    �                                         �    �                     S                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     '                    �    �                     \                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     0                    �    �                     e                    �    �                     �                    �    �                     �                    �    �                                         �    �                     9                    �    �                     n                    �    �                     �                    �    �                     �                    �    �                                         �    �                     B                    �    �                     w                    �    �                      �                     �    �                      �                     �    �                     �                    �    �                     �                    �    �                                         �    �                     0                    �    �                     S                    �    �                     v                    �    �                     �                    �    �                     �                    �    �                      �                     �    �                      �                     �    �                                           �    �                      7                     �    �                      g                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      '                     �    �                      W                     5�_�  3  5          4   7       ����                                                                                                                                                                                                                                                                                                                7           �          6          V       f�     �   5   6   �   �           -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  o      �   5   �       �       -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   6       �       5             j             �    5                                          5�_�  4  6          5   6       ����                                                                                                                                                                                                                                                                                                                6           �          5          V       f�     �   4   5   �   �       -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  n      �   4   �       �       -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   5       �       4              f      �      5�_�  5  7          6   5       ����                                                                                                                                                                                                                                                                                                                5           �          4          V       f�     �   3   4   �   �       -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  m      �   3   �       �       -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   4       �       3       �      f      �      �    4                     �                    �    5                                         �    6                     H                    �    7                     s                    �    8                     �                    �    9                     �                    �    :                     �                    �    ;                                         �    <                     J                    �    =                     u                    �    >                     �                    �    ?                     �                    �    @                     �                    �    A                     #                    �    B                     O                    �    C                     {                    �    D                     �                    �    E                     �                    �    F                     �                    �    G                     +                    �    H                     W                    �    I                     �                    �    J                     �                    �    K                     �                    �    L                     	                    �    M                     3	                    �    N                     _	                    �    O                     �	                    �    P                     �	                    �    Q                     �	                    �    R                     
                    �    S                     ;
                    �    T                     g
                    �    U                     �
                    �    V                     �
                    �    W                     �
                    �    X                                         �    Y                     C                    �    Z                     o                    �    [                     �                    �    \                     �                    �    ]                     �                    �    ^                                         �    _                     K                    �    `                     w                    �    a                     �                    �    b                     �                    �    c                     �                    �    d                     '                    �    e                     S                    �    f                                         �    g                     �                    �    h                     �                    �    i                                         �    j                     /                    �    k                     [                    �    l                     �                    �    m                     �                    �    n                     �                    �    o                                         �    p                     7                    �    q                     c                    �    r                     �                    �    s                     �                    �    t                     �                    �    u                                         �    w                     (                    �    x                     K                    �    y                     �                    �    z                     �                    �    {                     �                    �    |                     +                    �    }                     c                    �    ~                     �                    �                         �                    �    �                                         �    �                     C                    �    �                     {                    �    �                     �                    �    �                     �                    �    �                     &                    �    �                     _                    �    �                     �                    �    �                     �                    �    �                     
                    �    �                     C                    �    �                     |                    �    �                     �                    �    �                     �                    �    �                     '                    �    �                     `                    �    �                     �                    �    �                     �                    �    �                                         �    �                     D                    �    �                     }                    �    �                     �                    �    �                     �                    �    �                     (                    �    �                     a                    �    �                     �                    �    �                     �                    �    �                                         �    �                     E                    �    �                     ~                    �    �                     �                    �    �                     �                    �    �                     )                    �    �                     b                    �    �                     �                    �    �                     �                    �    �                                         �    �                     F                    �    �                                         �    �                     �                    �    �                     �                    �    �                     *                    �    �                     c                    �    �                     �                    �    �                     �                    �    �                                         �    �                     G                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     +                    �    �                     d                    �    �                     �                    �    �                     �                    �    �                                         �    �                     H                    �    �                      �                     �    �                      �                     �    �                     �                    �    �                     �                    �    �                     �                    �    �                                         �    �                     @                    �    �                     g                    �    �                     �                    �    �                     �                    �    �                      �                     �    �                      �                     �    �                                            �    �                      @                      �    �                      t                      �    �                      �                      �    �                      �                      �    �                      !                     �    �                      D!                     �    �                      x!                     5�_�  6  8          7   4       ����                                                                                                                                                                                                                                                                                                                4           �          3          V       f�     �   2   3   �   �       -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  l      �   2   �       �           -- Constants   #            type k_vector is record   .                K_0 : bit_vector(31 downto 0);   .                K_1 : bit_vector(31 downto 0);   .                K_2 : bit_vector(31 downto 0);   .                K_3 : bit_vector(31 downto 0);   .                K_4 : bit_vector(31 downto 0);   .                K_5 : bit_vector(31 downto 0);   .                K_6 : bit_vector(31 downto 0);   .                K_7 : bit_vector(31 downto 0);   .                K_8 : bit_vector(31 downto 0);   .                K_9 : bit_vector(31 downto 0);   /                K_10 : bit_vector(31 downto 0);   /                K_11 : bit_vector(31 downto 0);   /                K_12 : bit_vector(31 downto 0);   /                K_13 : bit_vector(31 downto 0);   /                K_14 : bit_vector(31 downto 0);   /                K_15 : bit_vector(31 downto 0);   /                K_16 : bit_vector(31 downto 0);   /                K_17 : bit_vector(31 downto 0);   /                K_18 : bit_vector(31 downto 0);   /                K_19 : bit_vector(31 downto 0);   /                K_20 : bit_vector(31 downto 0);   /                K_21 : bit_vector(31 downto 0);   /                K_22 : bit_vector(31 downto 0);   /                K_23 : bit_vector(31 downto 0);   /                K_24 : bit_vector(31 downto 0);   /                K_25 : bit_vector(31 downto 0);   /                K_26 : bit_vector(31 downto 0);   /                K_27 : bit_vector(31 downto 0);   /                K_28 : bit_vector(31 downto 0);   /                K_29 : bit_vector(31 downto 0);   /                K_30 : bit_vector(31 downto 0);   /                K_31 : bit_vector(31 downto 0);   /                K_32 : bit_vector(31 downto 0);   /                K_33 : bit_vector(31 downto 0);   /                K_34 : bit_vector(31 downto 0);   /                K_35 : bit_vector(31 downto 0);   /                K_36 : bit_vector(31 downto 0);   /                K_37 : bit_vector(31 downto 0);   /                K_38 : bit_vector(31 downto 0);   /                K_39 : bit_vector(31 downto 0);   /                K_40 : bit_vector(31 downto 0);   /                K_41 : bit_vector(31 downto 0);   /                K_42 : bit_vector(31 downto 0);   /                K_43 : bit_vector(31 downto 0);   /                K_44 : bit_vector(31 downto 0);   /                K_45 : bit_vector(31 downto 0);   /                K_46 : bit_vector(31 downto 0);   /                K_47 : bit_vector(31 downto 0);   /                K_48 : bit_vector(31 downto 0);   /                K_49 : bit_vector(31 downto 0);   /                K_50 : bit_vector(31 downto 0);   /                K_51 : bit_vector(31 downto 0);   /                K_52 : bit_vector(31 downto 0);   /                K_53 : bit_vector(31 downto 0);   /                K_54 : bit_vector(31 downto 0);   /                K_55 : bit_vector(31 downto 0);   /                K_56 : bit_vector(31 downto 0);   /                K_57 : bit_vector(31 downto 0);   /                K_58 : bit_vector(31 downto 0);   /                K_59 : bit_vector(31 downto 0);   /                K_60 : bit_vector(31 downto 0);   /                K_61 : bit_vector(31 downto 0);   /                K_62 : bit_vector(31 downto 0);   /                K_63 : bit_vector(31 downto 0);               end record;       &            constant K : k_vector := (   ;            K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   ;            K_1 => bit_vector(to_signed(32, 16#71374491#)),   ;            K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   ;            K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   ;            K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   ;            K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   ;            K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   ;            K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   ;            K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   ;            K_9 => bit_vector(to_signed(32, 16#12835b01#)),   <            K_10 => bit_vector(to_signed(32, 16#243185be#)),   <            K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   <            K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   <            K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   <            K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   <            K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   <            K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   <            K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   <            K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   <            K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   <            K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   <            K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   <            K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   <            K_23 => bit_vector(to_signed(32, 16#76f988da#)),   <            K_24 => bit_vector(to_signed(32, 16#983e5152#)),   <            K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   <            K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   <            K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   <            K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   <            K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   <            K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   <            K_31 => bit_vector(to_signed(32, 16#14292967#)),   <            K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   <            K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   <            K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   <            K_35 => bit_vector(to_signed(32, 16#53380d13#)),   <            K_36 => bit_vector(to_signed(32, 16#650a7354#)),   <            K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   <            K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   <            K_39 => bit_vector(to_signed(32, 16#92722c85#)),   <            K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   <            K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   <            K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   <            K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   <            K_44 => bit_vector(to_signed(32, 16#d192e819#)),   <            K_45 => bit_vector(to_signed(32, 16#d6990624#)),   <            K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   <            K_47 => bit_vector(to_signed(32, 16#106aa070#)),   <            K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   <            K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   <            K_50 => bit_vector(to_signed(32, 16#2748774c#)),   <            K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   <            K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   <            K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   <            K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   <            K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   <            K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   <            K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   <            K_58 => bit_vector(to_signed(32, 16#84c87814#)),   <            K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   <            K_60 => bit_vector(to_signed(32, 16#90befffa#)),   <            K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   <            K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   ;            K_63 => bit_vector(to_signed(32, 16#c67178f2#))   
        );               type h_vector is record   *            H_0 : bit_vector(31 downto 0);   *            H_1 : bit_vector(31 downto 0);   *            H_2 : bit_vector(31 downto 0);   *            H_3 : bit_vector(31 downto 0);   *            H_4 : bit_vector(31 downto 0);   *            H_5 : bit_vector(31 downto 0);   *            H_6 : bit_vector(31 downto 0);   *            H_7 : bit_vector(31 downto 0);           end record;       "        constant H : h_vector := (   7        H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   7        H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   7        H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   7        H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   7        H_4 => bit_vector(to_signed(32, 16#510e527f#)),   7        H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   7        H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   6        H_7 => bit_vector(to_signed(32, 16#5be0cd19#))       );5��   3       �       2       �      �      �      �    2                     �                    �    3                     �                    �    4                                         �    5                     I                    �    6                     x                    �    7                     �                    �    8                     �                    �    9                                         �    :                     4                    �    ;                     c                    �    <                     �                    �    =                     �                    �    >                     �                    �    ?                                          �    @                     P                    �    A                     �                    �    B                     �                    �    C                     �                    �    D                                         �    E                     @                    �    F                     p                    �    G                     �                    �    H                     �                    �    I                      	                    �    J                     0	                    �    K                     `	                    �    L                     �	                    �    M                     �	                    �    N                     �	                    �    O                      
                    �    P                     P
                    �    Q                     �
                    �    R                     �
                    �    S                     �
                    �    T                                         �    U                     @                    �    V                     p                    �    W                     �                    �    X                     �                    �    Y                                          �    Z                     0                    �    [                     `                    �    \                     �                    �    ]                     �                    �    ^                     �                    �    _                                          �    `                     P                    �    a                     �                    �    b                     �                    �    c                     �                    �    d                                         �    e                     @                    �    f                     p                    �    g                     �                    �    h                     �                    �    i                                          �    j                     0                    �    k                     `                    �    l                     �                    �    m                     �                    �    n                     �                    �    o                                          �    p                     P                    �    q                     �                    �    r                     �                    �    s                     �                    �    t                                         �    v                     )                    �    w                     P                    �    x                     �                    �    y                     �                    �    z                                         �    {                     @                    �    |                     |                    �    }                     �                    �    ~                     �                    �                         0                    �    �                     l                    �    �                     �                    �    �                     �                    �    �                     "                    �    �                     _                    �    �                     �                    �    �                     �                    �    �                                         �    �                     S                    �    �                     �                    �    �                     �                    �    �                     
                    �    �                     G                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     ;                    �    �                     x                    �    �                     �                    �    �                     �                    �    �                     /                    �    �                     l                    �    �                     �                    �    �                     �                    �    �                     #                    �    �                     `                    �    �                     �                    �    �                     �                    �    �                                         �    �                     T                    �    �                     �                    �    �                     �                    �    �                                         �    �                     H                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     <                    �    �                     y                    �    �                     �                    �    �                     �                    �    �                     0                    �    �                     m                    �    �                     �                    �    �                     �                    �    �                     $                    �    �                     a                    �    �                     �                    �    �                     �                    �    �                                         �    �                     U                    �    �                     �                    �    �                     �                    �    �                                          �    �                     I                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     !                    �    �                     2!                    �    �                     ]!                    �    �                     �!                    �    �                     �!                    �    �                     �!                    �    �                     	"                    �    �                     "                    �    �                     A"                    �    �                     y"                    �    �                     �"                    �    �                     �"                    �    �                     !#                    �    �                     Y#                    �    �                     �#                    �    �                     �#                    �    �                       $                     5�_�  7  9          8   3       ����                                                                                                                                                                                                                                                                                                                3           �          2          V       f�     �   1   2   �   �           -- Constants   #            type k_vector is record   .                K_0 : bit_vector(31 downto 0);   .                K_1 : bit_vector(31 downto 0);   .                K_2 : bit_vector(31 downto 0);   .                K_3 : bit_vector(31 downto 0);   .                K_4 : bit_vector(31 downto 0);   .                K_5 : bit_vector(31 downto 0);   .                K_6 : bit_vector(31 downto 0);   .                K_7 : bit_vector(31 downto 0);   .                K_8 : bit_vector(31 downto 0);   .                K_9 : bit_vector(31 downto 0);   /                K_10 : bit_vector(31 downto 0);   /                K_11 : bit_vector(31 downto 0);   /                K_12 : bit_vector(31 downto 0);   /                K_13 : bit_vector(31 downto 0);   /                K_14 : bit_vector(31 downto 0);   /                K_15 : bit_vector(31 downto 0);   /                K_16 : bit_vector(31 downto 0);   /                K_17 : bit_vector(31 downto 0);   /                K_18 : bit_vector(31 downto 0);   /                K_19 : bit_vector(31 downto 0);   /                K_20 : bit_vector(31 downto 0);   /                K_21 : bit_vector(31 downto 0);   /                K_22 : bit_vector(31 downto 0);   /                K_23 : bit_vector(31 downto 0);   /                K_24 : bit_vector(31 downto 0);   /                K_25 : bit_vector(31 downto 0);   /                K_26 : bit_vector(31 downto 0);   /                K_27 : bit_vector(31 downto 0);   /                K_28 : bit_vector(31 downto 0);   /                K_29 : bit_vector(31 downto 0);   /                K_30 : bit_vector(31 downto 0);   /                K_31 : bit_vector(31 downto 0);   /                K_32 : bit_vector(31 downto 0);   /                K_33 : bit_vector(31 downto 0);   /                K_34 : bit_vector(31 downto 0);   /                K_35 : bit_vector(31 downto 0);   /                K_36 : bit_vector(31 downto 0);   /                K_37 : bit_vector(31 downto 0);   /                K_38 : bit_vector(31 downto 0);   /                K_39 : bit_vector(31 downto 0);   /                K_40 : bit_vector(31 downto 0);   /                K_41 : bit_vector(31 downto 0);   /                K_42 : bit_vector(31 downto 0);   /                K_43 : bit_vector(31 downto 0);   /                K_44 : bit_vector(31 downto 0);   /                K_45 : bit_vector(31 downto 0);   /                K_46 : bit_vector(31 downto 0);   /                K_47 : bit_vector(31 downto 0);   /                K_48 : bit_vector(31 downto 0);   /                K_49 : bit_vector(31 downto 0);   /                K_50 : bit_vector(31 downto 0);   /                K_51 : bit_vector(31 downto 0);   /                K_52 : bit_vector(31 downto 0);   /                K_53 : bit_vector(31 downto 0);   /                K_54 : bit_vector(31 downto 0);   /                K_55 : bit_vector(31 downto 0);   /                K_56 : bit_vector(31 downto 0);   /                K_57 : bit_vector(31 downto 0);   /                K_58 : bit_vector(31 downto 0);   /                K_59 : bit_vector(31 downto 0);   /                K_60 : bit_vector(31 downto 0);   /                K_61 : bit_vector(31 downto 0);   /                K_62 : bit_vector(31 downto 0);   /                K_63 : bit_vector(31 downto 0);               end record;       &            constant K : k_vector := (   ;            K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   ;            K_1 => bit_vector(to_signed(32, 16#71374491#)),   ;            K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   ;            K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   ;            K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   ;            K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   ;            K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   ;            K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   ;            K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   ;            K_9 => bit_vector(to_signed(32, 16#12835b01#)),   <            K_10 => bit_vector(to_signed(32, 16#243185be#)),   <            K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   <            K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   <            K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   <            K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   <            K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   <            K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   <            K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   <            K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   <            K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   <            K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   <            K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   <            K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   <            K_23 => bit_vector(to_signed(32, 16#76f988da#)),   <            K_24 => bit_vector(to_signed(32, 16#983e5152#)),   <            K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   <            K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   <            K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   <            K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   <            K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   <            K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   <            K_31 => bit_vector(to_signed(32, 16#14292967#)),   <            K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   <            K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   <            K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   <            K_35 => bit_vector(to_signed(32, 16#53380d13#)),   <            K_36 => bit_vector(to_signed(32, 16#650a7354#)),   <            K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   <            K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   <            K_39 => bit_vector(to_signed(32, 16#92722c85#)),   <            K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   <            K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   <            K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   <            K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   <            K_44 => bit_vector(to_signed(32, 16#d192e819#)),   <            K_45 => bit_vector(to_signed(32, 16#d6990624#)),   <            K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   <            K_47 => bit_vector(to_signed(32, 16#106aa070#)),   <            K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   <            K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   <            K_50 => bit_vector(to_signed(32, 16#2748774c#)),   <            K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   <            K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   <            K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   <            K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   <            K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   <            K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   <            K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   <            K_58 => bit_vector(to_signed(32, 16#84c87814#)),   <            K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   <            K_60 => bit_vector(to_signed(32, 16#90befffa#)),   <            K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   <            K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   ;            K_63 => bit_vector(to_signed(32, 16#c67178f2#))   
        );               type h_vector is record   *            H_0 : bit_vector(31 downto 0);   *            H_1 : bit_vector(31 downto 0);   *            H_2 : bit_vector(31 downto 0);   *            H_3 : bit_vector(31 downto 0);   *            H_4 : bit_vector(31 downto 0);   *            H_5 : bit_vector(31 downto 0);   *            H_6 : bit_vector(31 downto 0);   *            H_7 : bit_vector(31 downto 0);           end record;       "        constant H : h_vector := (   7        H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   7        H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   7        H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   7        H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   7        H_4 => bit_vector(to_signed(32, 16#510e527f#)),   7        H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   7        H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   6        H_7 => bit_vector(to_signed(32, 16#5be0cd19#))       );�   �  k      �   1   �       �               -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   2       �       1       �      &      �      �    1                     �                    �    2                     �                    �    3                     �                    �    4                     �                    �    5                     (                    �    6                     S                    �    7                     ~                    �    8                     �                    �    9                     �                    �    :                     �                    �    ;                     *                    �    <                     U                    �    =                     �                    �    >                     �                    �    ?                     �                    �    @                                         �    A                     0                    �    B                     \                    �    C                     �                    �    D                     �                    �    E                     �                    �    F                                         �    G                     8                    �    H                     d                    �    I                     �                    �    J                     �                    �    K                     �                    �    L                     	                    �    M                     @	                    �    N                     l	                    �    O                     �	                    �    P                     �	                    �    Q                     �	                    �    R                     
                    �    S                     H
                    �    T                     t
                    �    U                     �
                    �    V                     �
                    �    W                     �
                    �    X                     $                    �    Y                     P                    �    Z                     |                    �    [                     �                    �    \                     �                    �    ]                                          �    ^                     ,                    �    _                     X                    �    `                     �                    �    a                     �                    �    b                     �                    �    c                                         �    d                     4                    �    e                     `                    �    f                     �                    �    g                     �                    �    h                     �                    �    i                                         �    j                     <                    �    k                     h                    �    l                     �                    �    m                     �                    �    n                     �                    �    o                                         �    p                     D                    �    q                     p                    �    r                     �                    �    s                     �                    �    u                     �                    �    v                                          �    w                     8                    �    x                     p                    �    y                     �                    �    z                     �                    �    {                                         �    |                     P                    �    }                     �                    �    ~                     �                    �                         �                    �    �                     0                    �    �                     i                    �    �                     �                    �    �                     �                    �    �                                         �    �                     M                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     1                    �    �                     j                    �    �                     �                    �    �                     �                    �    �                                         �    �                     N                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     2                    �    �                     k                    �    �                     �                    �    �                     �                    �    �                                         �    �                     O                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     3                    �    �                     l                    �    �                     �                    �    �                     �                    �    �                                         �    �                     P                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     4                    �    �                     m                    �    �                     �                    �    �                     �                    �    �                                         �    �                     Q                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     5                    �    �                     n                    �    �                     �                    �    �                     �                    �    �                                         �    �                     R                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     5                    �    �                     =                    �    �                     Y                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                                         �    �                     C                    �    �                     j                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     )                     �    �                     ]                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     -!                    �    �                      `!                     5�_�  8  :          9   2       ����                                                                                                                                                                                                                                                                                                                2           �          1          V       f�     �   0   1   �   �               -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  j      �   0   �       �           -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   1       �       0       �      �      l      �    0                     l                    5�_�  9  ;          :   1       ����                                                                                                                                                                                                                                                                                                                1           �          0          V       f�     �   /   0   �   �           -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  i      �   /   �       �           -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   0       �       /       l      �      '      5�_�  :  <          ;   0       ����                                                                                                                                                                                                                                                                                                                0           �          /          V       f�     �   .   /   �   �           -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  h      �   .   �       �           -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   /       �       .       '      �            �    /                     -                    �    0                     I                    �    1                     p                    �    2                     �                    �    3                     �                    �    4                     �                    �    5                                         �    6                     3                    �    7                     Z                    �    8                     �                    �    9                     �                    �    :                     �                    �    ;                     �                    �    <                                         �    =                     G                    �    >                     o                    �    ?                     �                    �    @                     �                    �    A                     �                    �    B                                         �    C                     7                    �    D                     _                    �    E                     �                    �    F                     �                    �    G                     �                    �    H                     �                    �    I                     '                    �    J                     O                    �    K                     w                    �    L                     �                    �    M                     �                    �    N                     �                    �    O                     	                    �    P                     ?	                    �    Q                     g	                    �    R                     �	                    �    S                     �	                    �    T                     �	                    �    U                     
                    �    V                     /
                    �    W                     W
                    �    X                     
                    �    Y                     �
                    �    Z                     �
                    �    [                     �
                    �    \                                         �    ]                     G                    �    ^                     o                    �    _                     �                    �    `                     �                    �    a                     �                    �    b                                         �    c                     7                    �    d                     _                    �    e                     �                    �    f                     �                    �    g                     �                    �    h                     �                    �    i                     '                    �    j                     O                    �    k                     w                    �    l                     �                    �    m                     �                    �    n                     �                    �    o                                         �    p                     ?                    �    r                     P                    �    s                     o                    �    t                     �                    �    u                     �                    �    v                                         �    w                     ?                    �    x                     s                    �    y                     �                    �    z                     �                    �    {                                         �    |                     C                    �    }                     w                    �    ~                     �                    �                         �                    �    �                                         �    �                     K                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                                         �    �                     T                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     (                    �    �                     ]                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     1                    �    �                     f                    �    �                     �                    �    �                     �                    �    �                                         �    �                     :                    �    �                     o                    �    �                     �                    �    �                     �                    �    �                                         �    �                     C                    �    �                     x                    �    �                     �                    �    �                     �                    �    �                                         �    �                     L                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                                          �    �                     U                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     )                    �    �                     ^                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     2                    �    �                     g                    �    �                     �                    �    �                     �                    �    �                                         �    �                     ;                    �    �                     p                    �    �                      �                     �    �                      �                     �    �                     �                    �    �                     �                    �    �                                         �    �                     )                    �    �                     L                    �    �                     o                    �    �                     �                    �    �                     �                    �    �                      �                     �    �                      �                     �    �                                            �    �                      0                     �    �                      `                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                                            �    �                      P                     5�_�  ;  =          <   /       ����                                                                                                                                                                                                                                                                                                                /           �          .          V       f�     �   -   .   �   �           -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  g      �   -   �       �       -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   .       �       -             j      �      �    -                     �                    �    .                                           �    /                     '                    �    0                     J                    �    1                     m                    �    2                     �                    �    3                     �                    �    4                     �                    �    5                     �                    �    6                                         �    7                     ?                    �    8                     b                    �    9                     �                    �    :                     �                    �    ;                     �                    �    <                     �                    �    =                                         �    >                     9                    �    ?                     ]                    �    @                     �                    �    A                     �                    �    B                     �                    �    C                     �                    �    D                                         �    E                     5                    �    F                     Y                    �    G                     }                    �    H                     �                    �    I                     �                    �    J                     �                    �    K                                         �    L                     1                    �    M                     U                    �    N                     y                    �    O                     �                    �    P                     �                    �    Q                     �                    �    R                     		                    �    S                     -	                    �    T                     Q	                    �    U                     u	                    �    V                     �	                    �    W                     �	                    �    X                     �	                    �    Y                     
                    �    Z                     )
                    �    [                     M
                    �    \                     q
                    �    ]                     �
                    �    ^                     �
                    �    _                     �
                    �    `                                         �    a                     %                    �    b                     I                    �    c                     m                    �    d                     �                    �    e                     �                    �    f                     �                    �    g                     �                    �    h                     !                    �    i                     E                    �    j                     i                    �    k                     �                    �    l                     �                    �    m                     �                    �    n                     �                    �    o                                           �    q                      *                     �    r                      E                     �    s                      u                     �    t                      �                     �    u                      �                     �    v                                           �    w                      5                     �    x                      e                     �    y                      �                     �    z                      �                     �    {                      �                     �    |                      %                     �    }                      V                     �    ~                      �                     �                          �                     �    �                      �                     �    �                                           �    �                      K                     �    �                      |                     �    �                      �                     �    �                      �                     �    �                                           �    �                      @                     �    �                      q                     �    �                      �                     �    �                      �                     �    �                                           �    �                      5                     �    �                      f                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      *                     �    �                      [                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                                           �    �                      P                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                                           �    �                      E                     �    �                      v                     �    �                      �                     �    �                      �                     �    �                      	                     �    �                      :                     �    �                      k                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      /                     �    �                      `                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      $                     �    �                      U                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                                           �    �                      J                     5�_�  <  >          =   .       ����                                                                                                                                                                                                                                                                                                                .           �          -          V       f�     �   ,   -   �   �       -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  f      �   ,   �       �   -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   -       �       ,       �      Z      �      �    ,                      �                     5�_�  =  ?          >   -       ����                                                                                                                                                                                                                                                                                                                -           �          ,          V       f�     �   +   ,   �   �   -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  e      �   +   �       �   -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   ,       �       +       �      V      �      5�_�  >  @          ?   ,       ����                                                                                                                                                                                                                                                                                                                ,           �          +          V       f�     �   *   +   �   �   -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  d      �   *   �       �   -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   +       �       *       �      V      �      5�_�  ?  A          @   +       ����                                                                                                                                                                                                                                                                                                                +           �          *          V       f�     �   )   *   �   �   -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  c      �   )   �       �   -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   *       �       )       �      V      �      �    *                      �                     �    +                     �                    �    ,                                         �    -                     A                    �    .                     h                    �    /                     �                    �    0                     �                    �    1                     �                    �    2                                         �    3                     +                    �    4                     R                    �    5                     y                    �    6                     �                    �    7                     �                    �    8                     �                    �    9                                         �    :                     A                    �    ;                     i                    �    <                     �                    �    =                     �                    �    >                     �                    �    ?                     	                    �    @                     1                    �    A                     Y                    �    B                     �                    �    C                     �                    �    D                     �                    �    E                     �                    �    F                     !                    �    G                     I                    �    H                     q                    �    I                     �                    �    J                     �                    �    K                     �                    �    L                     	                    �    M                     9	                    �    N                     a	                    �    O                     �	                    �    P                     �	                    �    Q                     �	                    �    R                     
                    �    S                     )
                    �    T                     Q
                    �    U                     y
                    �    V                     �
                    �    W                     �
                    �    X                     �
                    �    Y                                         �    Z                     A                    �    [                     i                    �    \                     �                    �    ]                     �                    �    ^                     �                    �    _                     	                    �    `                     1                    �    a                     Y                    �    b                     �                    �    c                     �                    �    d                     �                    �    e                     �                    �    f                     !                    �    g                     I                    �    h                     q                    �    i                     �                    �    j                     �                    �    k                      �                     �    m                      �                     �    n                                           �    o                      M                     �    p                      �                     �    q                      �                     �    r                      �                     �    s                                           �    t                      Q                     �    u                      �                     �    v                      �                     �    w                      �                     �    x                      !                     �    y                      V                     �    z                      �                     �    {                      �                     �    |                      �                     �    }                      *                     �    ~                      _                     �                          �                     �    �                      �                     �    �                      �                     �    �                      3                     �    �                      h                     �    �                      �                     �    �                      �                     �    �                                           �    �                      <                     �    �                      q                     �    �                      �                     �    �                      �                     �    �                                           �    �                      E                     �    �                      z                     �    �                      �                     �    �                      �                     �    �                                           �    �                      N                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      "                     �    �                      W                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      +                     �    �                      `                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      4                     �    �                      i                     �    �                      �                     �    �                      �                     �    �                                           �    �                      =                     �    �                      r                     �    �                      �                     �    �                      �                     �    �                                           �    �                      F                     �    �                      {                     �    �                      �                     �    �                      �                     �    �                                           5�_�  @  B          A   *       ����                                                                                                                                                                                                                                                                                                                *           �          )          V       f�     �   (   )   �   �   -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  b      �   (   �       �       -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   )       �       (       �      b      �      �    (                      �                     �    )                     �                    �    *                     �                    �    +                                         �    ,                     J                    �    -                     u                    �    .                     �                    �    /                     �                    �    0                     �                    �    1                     !                    �    2                     L                    �    3                     w                    �    4                     �                    �    5                     �                    �    6                     �                    �    7                     &                    �    8                     R                    �    9                     ~                    �    :                     �                    �    ;                     �                    �    <                                         �    =                     .                    �    >                     Z                    �    ?                     �                    �    @                     �                    �    A                     �                    �    B                     
                    �    C                     6                    �    D                     b                    �    E                     �                    �    F                     �                    �    G                     �                    �    H                     	                    �    I                     >	                    �    J                     j	                    �    K                     �	                    �    L                     �	                    �    M                     �	                    �    N                     
                    �    O                     F
                    �    P                     r
                    �    Q                     �
                    �    R                     �
                    �    S                     �
                    �    T                     "                    �    U                     N                    �    V                     z                    �    W                     �                    �    X                     �                    �    Y                     �                    �    Z                     *                    �    [                     V                    �    \                     �                    �    ]                     �                    �    ^                     �                    �    _                                         �    `                     2                    �    a                     ^                    �    b                     �                    �    c                     �                    �    d                     �                    �    e                                         �    f                     :                    �    g                     f                    �    h                     �                    �    i                     �                    �    j                     �                    �    l                     �                    �    m                     "                    �    n                     Z                    �    o                     �                    �    p                     �                    �    q                                         �    r                     :                    �    s                     r                    �    t                     �                    �    u                     �                    �    v                                         �    w                     R                    �    x                     �                    �    y                     �                    �    z                     �                    �    {                     6                    �    |                     o                    �    }                     �                    �    ~                     �                    �                                             �    �                     S                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     7                    �    �                     p                    �    �                     �                    �    �                     �                    �    �                                         �    �                     T                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     8                    �    �                     q                    �    �                     �                    �    �                     �                    �    �                                         �    �                     U                    �    �                     �                    �    �                     �                    �    �                                          �    �                     9                    �    �                     r                    �    �                     �                    �    �                     �                    �    �                                         �    �                     V                    �    �                     �                    �    �                     �                    �    �                                         �    �                     :                    �    �                     s                    �    �                     �                    �    �                     �                    �    �                                         �    �                     W                    �    �                     �                    �    �                     �                    �    �                                         �    �                     ;                    �    �                     t                    �    �                     �                    �    �                     �                    �    �                                         �    �                      W                     �    �                      _                     �    �                     {                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                                         �    �                     >                    �    �                     e                    �    �                     �                    �    �                      �                     �    �                      �                     �    �                      �                     �    �                                           �    �                      K                     �    �                                           �    �                      �                     �    �                      �                     �    �                                            �    �                      O                      5�_�  A  C          B   )       ����                                                                                                                                                                                                                                                                                                                )           �          (          V       f�     �   '   (   �   �       -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  a      �   '   �       �           -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   (       �       '       �      �      �      �    '                     �                    �    (                     �                    �    )                     �                    �    *                                         �    +                     +                    �    ,                     R                    �    -                     y                    �    .                     �                    �    /                     �                    �    0                     �                    �    1                                         �    2                     <                    �    3                     c                    �    4                     �                    �    5                     �                    �    6                     �                    �    7                                         �    8                     +                    �    9                     S                    �    :                     {                    �    ;                     �                    �    <                     �                    �    =                     �                    �    >                                         �    ?                     C                    �    @                     k                    �    A                     �                    �    B                     �                    �    C                     �                    �    D                                         �    E                     3                    �    F                     [                    �    G                     �                    �    H                     �                    �    I                     �                    �    J                     �                    �    K                     #	                    �    L                     K	                    �    M                     s	                    �    N                     �	                    �    O                     �	                    �    P                     �	                    �    Q                     
                    �    R                     ;
                    �    S                     c
                    �    T                     �
                    �    U                     �
                    �    V                     �
                    �    W                                         �    X                     +                    �    Y                     S                    �    Z                     {                    �    [                     �                    �    \                     �                    �    ]                     �                    �    ^                                         �    _                     C                    �    `                     k                    �    a                     �                    �    b                     �                    �    c                     �                    �    d                                         �    e                     3                    �    f                     [                    �    g                     �                    �    h                     �                    �    i                     �                    �    k                     �                    �    l                                         �    m                     7                    �    n                     k                    �    o                     �                    �    p                     �                    �    q                                         �    r                     ;                    �    s                     o                    �    t                     �                    �    u                     �                    �    v                                         �    w                     @                    �    x                     u                    �    y                     �                    �    z                     �                    �    {                                         �    |                     I                    �    }                     ~                    �    ~                     �                    �                         �                    �    �                                         �    �                     R                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     &                    �    �                     [                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     /                    �    �                     d                    �    �                     �                    �    �                     �                    �    �                                         �    �                     8                    �    �                     m                    �    �                     �                    �    �                     �                    �    �                                         �    �                     A                    �    �                     v                    �    �                     �                    �    �                     �                    �    �                                         �    �                     J                    �    �                                         �    �                     �                    �    �                     �                    �    �                                         �    �                     S                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     '                    �    �                     \                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     0                    �    �                     e                    �    �                     �                    �    �                     �                    �    �                                         �    �                      8                     �    �                      <                     �    �                     T                    �    �                     w                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                                         �    �                     &                    �    �                     I                    �    �                      l                     �    �                      y                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      $                     �    �                      T                     �    �                      �                     �    �                      �                     �    �                      �                     5�_�  B  D          C   (       ����                                                                                                                                                                                                                                                                                                                (           �          '          V       f�     �   &   '   �   �           -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  `      �   &   �       �       -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   '       �       &       �      j            �    &                                         5�_�  C  E          D   '       ����                                                                                                                                                                                                                                                                                                                )           �          (          V       f�     �   �   �   �   �       -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   &   �      �   '   �       �       -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   &       �       '             f      �      5�_�  D  F          E   (       ����                                                                                                                                                                                                                                                                                                                *           �          )          V       f�     �   �   �   �   �       -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   '   �      �   (   �       �       -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   '       �       (       �      f      �      �    )                     �                    �    *                     �                    �    +                                         �    ,                     J                    �    -                     u                    �    .                     �                    �    /                     �                    �    0                     �                    �    1                     !                    �    2                     L                    �    3                     w                    �    4                     �                    �    5                     �                    �    6                     �                    �    7                     &                    �    8                     R                    �    9                     ~                    �    :                     �                    �    ;                     �                    �    <                                         �    =                     .                    �    >                     Z                    �    ?                     �                    �    @                     �                    �    A                     �                    �    B                     
                    �    C                     6                    �    D                     b                    �    E                     �                    �    F                     �                    �    G                     �                    �    H                     	                    �    I                     >	                    �    J                     j	                    �    K                     �	                    �    L                     �	                    �    M                     �	                    �    N                     
                    �    O                     F
                    �    P                     r
                    �    Q                     �
                    �    R                     �
                    �    S                     �
                    �    T                     "                    �    U                     N                    �    V                     z                    �    W                     �                    �    X                     �                    �    Y                     �                    �    Z                     *                    �    [                     V                    �    \                     �                    �    ]                     �                    �    ^                     �                    �    _                                         �    `                     2                    �    a                     ^                    �    b                     �                    �    c                     �                    �    d                     �                    �    e                                         �    f                     :                    �    g                     f                    �    h                     �                    �    i                     �                    �    j                     �                    �    l                     �                    �    m                     "                    �    n                     Z                    �    o                     �                    �    p                     �                    �    q                                         �    r                     :                    �    s                     r                    �    t                     �                    �    u                     �                    �    v                                         �    w                     R                    �    x                     �                    �    y                     �                    �    z                     �                    �    {                     6                    �    |                     o                    �    }                     �                    �    ~                     �                    �                                             �    �                     S                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     7                    �    �                     p                    �    �                     �                    �    �                     �                    �    �                                         �    �                     T                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     8                    �    �                     q                    �    �                     �                    �    �                     �                    �    �                                         �    �                     U                    �    �                     �                    �    �                     �                    �    �                                          �    �                     9                    �    �                     r                    �    �                     �                    �    �                     �                    �    �                                         �    �                     V                    �    �                     �                    �    �                     �                    �    �                                         �    �                     :                    �    �                     s                    �    �                     �                    �    �                     �                    �    �                                         �    �                     W                    �    �                     �                    �    �                     �                    �    �                                         �    �                     ;                    �    �                     t                    �    �                     �                    �    �                     �                    �    �                                         �    �                      W                     �    �                      _                     �    �                     {                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                                         �    �                     >                    �    �                     e                    �    �                     �                    �    �                      �                     �    �                      �                     �    �                      �                     �    �                                           �    �                      K                     �    �                                           �    �                      �                     �    �                      �                     �    �                                            �    �                      O                      5�_�  E  G          F   )       ����                                                                                                                                                                                                                                                                                                                +           �          *          V       f�     �   �   �   �   �       -- Constants           type k_vector is record   *            K_0 : bit_vector(31 downto 0);   *            K_1 : bit_vector(31 downto 0);   *            K_2 : bit_vector(31 downto 0);   *            K_3 : bit_vector(31 downto 0);   *            K_4 : bit_vector(31 downto 0);   *            K_5 : bit_vector(31 downto 0);   *            K_6 : bit_vector(31 downto 0);   *            K_7 : bit_vector(31 downto 0);   *            K_8 : bit_vector(31 downto 0);   *            K_9 : bit_vector(31 downto 0);   +            K_10 : bit_vector(31 downto 0);   +            K_11 : bit_vector(31 downto 0);   +            K_12 : bit_vector(31 downto 0);   +            K_13 : bit_vector(31 downto 0);   +            K_14 : bit_vector(31 downto 0);   +            K_15 : bit_vector(31 downto 0);   +            K_16 : bit_vector(31 downto 0);   +            K_17 : bit_vector(31 downto 0);   +            K_18 : bit_vector(31 downto 0);   +            K_19 : bit_vector(31 downto 0);   +            K_20 : bit_vector(31 downto 0);   +            K_21 : bit_vector(31 downto 0);   +            K_22 : bit_vector(31 downto 0);   +            K_23 : bit_vector(31 downto 0);   +            K_24 : bit_vector(31 downto 0);   +            K_25 : bit_vector(31 downto 0);   +            K_26 : bit_vector(31 downto 0);   +            K_27 : bit_vector(31 downto 0);   +            K_28 : bit_vector(31 downto 0);   +            K_29 : bit_vector(31 downto 0);   +            K_30 : bit_vector(31 downto 0);   +            K_31 : bit_vector(31 downto 0);   +            K_32 : bit_vector(31 downto 0);   +            K_33 : bit_vector(31 downto 0);   +            K_34 : bit_vector(31 downto 0);   +            K_35 : bit_vector(31 downto 0);   +            K_36 : bit_vector(31 downto 0);   +            K_37 : bit_vector(31 downto 0);   +            K_38 : bit_vector(31 downto 0);   +            K_39 : bit_vector(31 downto 0);   +            K_40 : bit_vector(31 downto 0);   +            K_41 : bit_vector(31 downto 0);   +            K_42 : bit_vector(31 downto 0);   +            K_43 : bit_vector(31 downto 0);   +            K_44 : bit_vector(31 downto 0);   +            K_45 : bit_vector(31 downto 0);   +            K_46 : bit_vector(31 downto 0);   +            K_47 : bit_vector(31 downto 0);   +            K_48 : bit_vector(31 downto 0);   +            K_49 : bit_vector(31 downto 0);   +            K_50 : bit_vector(31 downto 0);   +            K_51 : bit_vector(31 downto 0);   +            K_52 : bit_vector(31 downto 0);   +            K_53 : bit_vector(31 downto 0);   +            K_54 : bit_vector(31 downto 0);   +            K_55 : bit_vector(31 downto 0);   +            K_56 : bit_vector(31 downto 0);   +            K_57 : bit_vector(31 downto 0);   +            K_58 : bit_vector(31 downto 0);   +            K_59 : bit_vector(31 downto 0);   +            K_60 : bit_vector(31 downto 0);   +            K_61 : bit_vector(31 downto 0);   +            K_62 : bit_vector(31 downto 0);   +            K_63 : bit_vector(31 downto 0);           end record;       "        constant K : k_vector := (   7        K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   7        K_1 => bit_vector(to_signed(32, 16#71374491#)),   7        K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   7        K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   7        K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   7        K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   7        K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   7        K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   7        K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   7        K_9 => bit_vector(to_signed(32, 16#12835b01#)),   8        K_10 => bit_vector(to_signed(32, 16#243185be#)),   8        K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   8        K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   8        K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   8        K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   8        K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   8        K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   8        K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   8        K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   8        K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   8        K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   8        K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   8        K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   8        K_23 => bit_vector(to_signed(32, 16#76f988da#)),   8        K_24 => bit_vector(to_signed(32, 16#983e5152#)),   8        K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   8        K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   8        K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   8        K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   8        K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   8        K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   8        K_31 => bit_vector(to_signed(32, 16#14292967#)),   8        K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   8        K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   8        K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   8        K_35 => bit_vector(to_signed(32, 16#53380d13#)),   8        K_36 => bit_vector(to_signed(32, 16#650a7354#)),   8        K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   8        K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   8        K_39 => bit_vector(to_signed(32, 16#92722c85#)),   8        K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   8        K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   8        K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   8        K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   8        K_44 => bit_vector(to_signed(32, 16#d192e819#)),   8        K_45 => bit_vector(to_signed(32, 16#d6990624#)),   8        K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   8        K_47 => bit_vector(to_signed(32, 16#106aa070#)),   8        K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   8        K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   8        K_50 => bit_vector(to_signed(32, 16#2748774c#)),   8        K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   8        K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   8        K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   8        K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   8        K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   8        K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   8        K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   8        K_58 => bit_vector(to_signed(32, 16#84c87814#)),   8        K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   8        K_60 => bit_vector(to_signed(32, 16#90befffa#)),   8        K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   8        K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   7        K_63 => bit_vector(to_signed(32, 16#c67178f2#))       );           type h_vector is record   &        H_0 : bit_vector(31 downto 0);   &        H_1 : bit_vector(31 downto 0);   &        H_2 : bit_vector(31 downto 0);   &        H_3 : bit_vector(31 downto 0);   &        H_4 : bit_vector(31 downto 0);   &        H_5 : bit_vector(31 downto 0);   &        H_6 : bit_vector(31 downto 0);   &        H_7 : bit_vector(31 downto 0);       end record;           constant H : h_vector := (   3    H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   3    H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   3    H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   3    H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   3    H_4 => bit_vector(to_signed(32, 16#510e527f#)),   3    H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   3    H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   2    H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   (   �      �   )   �       �           -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   (       �       )       �      �      �      �    )                     �                    �    *                     �                    �    +                     �                    �    ,                     "                    �    -                     I                    �    .                     p                    �    /                     �                    �    0                     �                    �    1                     �                    �    2                                         �    3                     3                    �    4                     Z                    �    5                     �                    �    6                     �                    �    7                     �                    �    8                     �                    �    9                     !                    �    :                     I                    �    ;                     q                    �    <                     �                    �    =                     �                    �    >                     �                    �    ?                                         �    @                     9                    �    A                     a                    �    B                     �                    �    C                     �                    �    D                     �                    �    E                                         �    F                     )                    �    G                     Q                    �    H                     y                    �    I                     �                    �    J                     �                    �    K                     �                    �    L                     	                    �    M                     A	                    �    N                     i	                    �    O                     �	                    �    P                     �	                    �    Q                     �	                    �    R                     	
                    �    S                     1
                    �    T                     Y
                    �    U                     �
                    �    V                     �
                    �    W                     �
                    �    X                     �
                    �    Y                     !                    �    Z                     I                    �    [                     q                    �    \                     �                    �    ]                     �                    �    ^                     �                    �    _                                         �    `                     9                    �    a                     a                    �    b                     �                    �    c                     �                    �    d                     �                    �    e                                         �    f                     )                    �    g                     Q                    �    h                     y                    �    i                     �                    �    j                     �                    �    k                     �                    �    m                                         �    n                     !                    �    o                     U                    �    p                     �                    �    q                     �                    �    r                     �                    �    s                     %                    �    t                     Y                    �    u                     �                    �    v                     �                    �    w                     �                    �    x                     )                    �    y                     ^                    �    z                     �                    �    {                     �                    �    |                     �                    �    }                     2                    �    ~                     g                    �                         �                    �    �                     �                    �    �                                         �    �                     ;                    �    �                     p                    �    �                     �                    �    �                     �                    �    �                                         �    �                     D                    �    �                     y                    �    �                     �                    �    �                     �                    �    �                                         �    �                     M                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     !                    �    �                     V                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     *                    �    �                     _                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     3                    �    �                     h                    �    �                     �                    �    �                     �                    �    �                                         �    �                     <                    �    �                     q                    �    �                     �                    �    �                     �                    �    �                                         �    �                     E                    �    �                     z                    �    �                     �                    �    �                     �                    �    �                                         �    �                     N                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     "                    �    �                      V                     �    �                      Z                     �    �                     r                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     !                    �    �                     D                    �    �                     g                    �    �                      �                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                                           �    �                      B                     �    �                      r                     �    �                      �                     �    �                      �                     �    �                                           5�_�  F  H          G   *       ����                                                                                                                                                                                                                                                                                                                ,           �          +          V       f�     �   �   �   �   �           -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   )   �      �   *   �       �       -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   )       �       *       �      j      �      �    *                     �                    �    +                      �                     �    ,                                         �    -                     &                    �    .                     I                    �    /                     l                    �    0                     �                    �    1                     �                    �    2                     �                    �    3                     �                    �    4                                         �    5                     >                    �    6                     a                    �    7                     �                    �    8                     �                    �    9                     �                    �    :                     �                    �    ;                                         �    <                     9                    �    =                     ]                    �    >                     �                    �    ?                     �                    �    @                     �                    �    A                     �                    �    B                                         �    C                     5                    �    D                     Y                    �    E                     }                    �    F                     �                    �    G                     �                    �    H                     �                    �    I                                         �    J                     1                    �    K                     U                    �    L                     y                    �    M                     �                    �    N                     �                    �    O                     �                    �    P                     		                    �    Q                     -	                    �    R                     Q	                    �    S                     u	                    �    T                     �	                    �    U                     �	                    �    V                     �	                    �    W                     
                    �    X                     )
                    �    Y                     M
                    �    Z                     q
                    �    [                     �
                    �    \                     �
                    �    ]                     �
                    �    ^                                         �    _                     %                    �    `                     I                    �    a                     m                    �    b                     �                    �    c                     �                    �    d                     �                    �    e                     �                    �    f                     !                    �    g                     E                    �    h                     i                    �    i                     �                    �    j                     �                    �    k                     �                    �    l                      �                     �    n                                           �    o                      !                     �    p                      Q                     �    q                      �                     �    r                      �                     �    s                      �                     �    t                                           �    u                      A                     �    v                      q                     �    w                      �                     �    x                      �                     �    y                                           �    z                      2                     �    {                      c                     �    |                      �                     �    }                      �                     �    ~                      �                     �                          '                     �    �                      X                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                                           �    �                      M                     �    �                      ~                     �    �                      �                     �    �                      �                     �    �                                           �    �                      B                     �    �                      s                     �    �                      �                     �    �                      �                     �    �                                           �    �                      7                     �    �                      h                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      ,                     �    �                      ]                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      !                     �    �                      R                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                                           �    �                      G                     �    �                      x                     �    �                      �                     �    �                      �                     �    �                                           �    �                      <                     �    �                      m                     �    �                      �                     �    �                      �                     �    �                                            �    �                      1                     �    �                      b                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      &                     5�_�  G  I          H   +       ����                                                                                                                                                                                                                                                                                                                -           �          ,          V       f�     �   �   �   �   �       -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   *   �      �   +   �       �   -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   *       �       +       �      Z      �      �    +                      �                     5�_�  H  J          I   ,       ����                                                                                                                                                                                                                                                                                                                .           �          -          V       f�     �   �   �   �   �   -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   +   �      �   ,   �       �   -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   +       �       ,       �      V      �      5�_�  I  K          J   -       ����                                                                                                                                                                                                                                                                                                                /           �          .          V       f�     �   �   �   �   �   -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   ,   �      �   -   �       �   -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   ,       �       -       �      V      �      5�_�  J  L          K   .       ����                                                                                                                                                                                                                                                                                                                0           �          /          V       f�     �   �   �   �   �   -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   -   �      �   .   �       �   -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   -       �       .       �      V            �    /                      %                     �    0                     A                    �    1                     h                    �    2                     �                    �    3                     �                    �    4                     �                    �    5                                         �    6                     +                    �    7                     R                    �    8                     y                    �    9                     �                    �    :                     �                    �    ;                     �                    �    <                                         �    =                     ?                    �    >                     g                    �    ?                     �                    �    @                     �                    �    A                     �                    �    B                                         �    C                     /                    �    D                     W                    �    E                                         �    F                     �                    �    G                     �                    �    H                     �                    �    I                                         �    J                     G                    �    K                     o                    �    L                     �                    �    M                     �                    �    N                     �                    �    O                     	                    �    P                     7	                    �    Q                     _	                    �    R                     �	                    �    S                     �	                    �    T                     �	                    �    U                     �	                    �    V                     '
                    �    W                     O
                    �    X                     w
                    �    Y                     �
                    �    Z                     �
                    �    [                     �
                    �    \                                         �    ]                     ?                    �    ^                     g                    �    _                     �                    �    `                     �                    �    a                     �                    �    b                                         �    c                     /                    �    d                     W                    �    e                                         �    f                     �                    �    g                     �                    �    h                     �                    �    i                                         �    j                     G                    �    k                     o                    �    l                     �                    �    m                     �                    �    n                     �                    �    o                                         �    p                      7                     �    r                      H                     �    s                      g                     �    t                      �                     �    u                      �                     �    v                                           �    w                      7                     �    x                      k                     �    y                      �                     �    z                      �                     �    {                                           �    |                      ;                     �    }                      o                     �    ~                      �                     �                          �                     �    �                                           �    �                      C                     �    �                      x                     �    �                      �                     �    �                      �                     �    �                                           �    �                      L                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                                            �    �                      U                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      )                     �    �                      ^                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      2                     �    �                      g                     �    �                      �                     �    �                      �                     �    �                                           �    �                      ;                     �    �                      p                     �    �                      �                     �    �                      �                     �    �                                           �    �                      D                     �    �                      y                     �    �                      �                     �    �                      �                     �    �                                           �    �                      M                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      !                     �    �                      V                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      *                     �    �                      _                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      3                     �    �                      h                     5�_�  K              L   /       ����                                                                                                                                                                                                                                                                                                                /                                            f�    �   -   .   �   �   -- Constants       type k_vector is record   &        K_0 : bit_vector(31 downto 0);   &        K_1 : bit_vector(31 downto 0);   &        K_2 : bit_vector(31 downto 0);   &        K_3 : bit_vector(31 downto 0);   &        K_4 : bit_vector(31 downto 0);   &        K_5 : bit_vector(31 downto 0);   &        K_6 : bit_vector(31 downto 0);   &        K_7 : bit_vector(31 downto 0);   &        K_8 : bit_vector(31 downto 0);   &        K_9 : bit_vector(31 downto 0);   '        K_10 : bit_vector(31 downto 0);   '        K_11 : bit_vector(31 downto 0);   '        K_12 : bit_vector(31 downto 0);   '        K_13 : bit_vector(31 downto 0);   '        K_14 : bit_vector(31 downto 0);   '        K_15 : bit_vector(31 downto 0);   '        K_16 : bit_vector(31 downto 0);   '        K_17 : bit_vector(31 downto 0);   '        K_18 : bit_vector(31 downto 0);   '        K_19 : bit_vector(31 downto 0);   '        K_20 : bit_vector(31 downto 0);   '        K_21 : bit_vector(31 downto 0);   '        K_22 : bit_vector(31 downto 0);   '        K_23 : bit_vector(31 downto 0);   '        K_24 : bit_vector(31 downto 0);   '        K_25 : bit_vector(31 downto 0);   '        K_26 : bit_vector(31 downto 0);   '        K_27 : bit_vector(31 downto 0);   '        K_28 : bit_vector(31 downto 0);   '        K_29 : bit_vector(31 downto 0);   '        K_30 : bit_vector(31 downto 0);   '        K_31 : bit_vector(31 downto 0);   '        K_32 : bit_vector(31 downto 0);   '        K_33 : bit_vector(31 downto 0);   '        K_34 : bit_vector(31 downto 0);   '        K_35 : bit_vector(31 downto 0);   '        K_36 : bit_vector(31 downto 0);   '        K_37 : bit_vector(31 downto 0);   '        K_38 : bit_vector(31 downto 0);   '        K_39 : bit_vector(31 downto 0);   '        K_40 : bit_vector(31 downto 0);   '        K_41 : bit_vector(31 downto 0);   '        K_42 : bit_vector(31 downto 0);   '        K_43 : bit_vector(31 downto 0);   '        K_44 : bit_vector(31 downto 0);   '        K_45 : bit_vector(31 downto 0);   '        K_46 : bit_vector(31 downto 0);   '        K_47 : bit_vector(31 downto 0);   '        K_48 : bit_vector(31 downto 0);   '        K_49 : bit_vector(31 downto 0);   '        K_50 : bit_vector(31 downto 0);   '        K_51 : bit_vector(31 downto 0);   '        K_52 : bit_vector(31 downto 0);   '        K_53 : bit_vector(31 downto 0);   '        K_54 : bit_vector(31 downto 0);   '        K_55 : bit_vector(31 downto 0);   '        K_56 : bit_vector(31 downto 0);   '        K_57 : bit_vector(31 downto 0);   '        K_58 : bit_vector(31 downto 0);   '        K_59 : bit_vector(31 downto 0);   '        K_60 : bit_vector(31 downto 0);   '        K_61 : bit_vector(31 downto 0);   '        K_62 : bit_vector(31 downto 0);   '        K_63 : bit_vector(31 downto 0);       end record;           constant K : k_vector := (   3    K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   3    K_1 => bit_vector(to_signed(32, 16#71374491#)),   3    K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   3    K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   3    K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   3    K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   3    K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   3    K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   3    K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   3    K_9 => bit_vector(to_signed(32, 16#12835b01#)),   4    K_10 => bit_vector(to_signed(32, 16#243185be#)),   4    K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   4    K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   4    K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   4    K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   4    K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   4    K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   4    K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   4    K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   4    K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   4    K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   4    K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   4    K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   4    K_23 => bit_vector(to_signed(32, 16#76f988da#)),   4    K_24 => bit_vector(to_signed(32, 16#983e5152#)),   4    K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   4    K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   4    K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   4    K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   4    K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   4    K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   4    K_31 => bit_vector(to_signed(32, 16#14292967#)),   4    K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   4    K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   4    K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   4    K_35 => bit_vector(to_signed(32, 16#53380d13#)),   4    K_36 => bit_vector(to_signed(32, 16#650a7354#)),   4    K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   4    K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   4    K_39 => bit_vector(to_signed(32, 16#92722c85#)),   4    K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   4    K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   4    K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   4    K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   4    K_44 => bit_vector(to_signed(32, 16#d192e819#)),   4    K_45 => bit_vector(to_signed(32, 16#d6990624#)),   4    K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   4    K_47 => bit_vector(to_signed(32, 16#106aa070#)),   4    K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   4    K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   4    K_50 => bit_vector(to_signed(32, 16#2748774c#)),   4    K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   4    K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   4    K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   4    K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   4    K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   4    K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   4    K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   4    K_58 => bit_vector(to_signed(32, 16#84c87814#)),   4    K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   4    K_60 => bit_vector(to_signed(32, 16#90befffa#)),   4    K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   4    K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   3    K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );�   �  g      �   -   �       �       -- Constants   type k_vector is record   "    K_0 : bit_vector(31 downto 0);   "    K_1 : bit_vector(31 downto 0);   "    K_2 : bit_vector(31 downto 0);   "    K_3 : bit_vector(31 downto 0);   "    K_4 : bit_vector(31 downto 0);   "    K_5 : bit_vector(31 downto 0);   "    K_6 : bit_vector(31 downto 0);   "    K_7 : bit_vector(31 downto 0);   "    K_8 : bit_vector(31 downto 0);   "    K_9 : bit_vector(31 downto 0);   #    K_10 : bit_vector(31 downto 0);   #    K_11 : bit_vector(31 downto 0);   #    K_12 : bit_vector(31 downto 0);   #    K_13 : bit_vector(31 downto 0);   #    K_14 : bit_vector(31 downto 0);   #    K_15 : bit_vector(31 downto 0);   #    K_16 : bit_vector(31 downto 0);   #    K_17 : bit_vector(31 downto 0);   #    K_18 : bit_vector(31 downto 0);   #    K_19 : bit_vector(31 downto 0);   #    K_20 : bit_vector(31 downto 0);   #    K_21 : bit_vector(31 downto 0);   #    K_22 : bit_vector(31 downto 0);   #    K_23 : bit_vector(31 downto 0);   #    K_24 : bit_vector(31 downto 0);   #    K_25 : bit_vector(31 downto 0);   #    K_26 : bit_vector(31 downto 0);   #    K_27 : bit_vector(31 downto 0);   #    K_28 : bit_vector(31 downto 0);   #    K_29 : bit_vector(31 downto 0);   #    K_30 : bit_vector(31 downto 0);   #    K_31 : bit_vector(31 downto 0);   #    K_32 : bit_vector(31 downto 0);   #    K_33 : bit_vector(31 downto 0);   #    K_34 : bit_vector(31 downto 0);   #    K_35 : bit_vector(31 downto 0);   #    K_36 : bit_vector(31 downto 0);   #    K_37 : bit_vector(31 downto 0);   #    K_38 : bit_vector(31 downto 0);   #    K_39 : bit_vector(31 downto 0);   #    K_40 : bit_vector(31 downto 0);   #    K_41 : bit_vector(31 downto 0);   #    K_42 : bit_vector(31 downto 0);   #    K_43 : bit_vector(31 downto 0);   #    K_44 : bit_vector(31 downto 0);   #    K_45 : bit_vector(31 downto 0);   #    K_46 : bit_vector(31 downto 0);   #    K_47 : bit_vector(31 downto 0);   #    K_48 : bit_vector(31 downto 0);   #    K_49 : bit_vector(31 downto 0);   #    K_50 : bit_vector(31 downto 0);   #    K_51 : bit_vector(31 downto 0);   #    K_52 : bit_vector(31 downto 0);   #    K_53 : bit_vector(31 downto 0);   #    K_54 : bit_vector(31 downto 0);   #    K_55 : bit_vector(31 downto 0);   #    K_56 : bit_vector(31 downto 0);   #    K_57 : bit_vector(31 downto 0);   #    K_58 : bit_vector(31 downto 0);   #    K_59 : bit_vector(31 downto 0);   #    K_60 : bit_vector(31 downto 0);   #    K_61 : bit_vector(31 downto 0);   #    K_62 : bit_vector(31 downto 0);   #    K_63 : bit_vector(31 downto 0);   end record;       constant K : k_vector := (   /K_0 => bit_vector(to_signed(32, 16#428a2f98#)),   /K_1 => bit_vector(to_signed(32, 16#71374491#)),   /K_2 => bit_vector(to_signed(32, 16#b5c0fbcf#)),   /K_3 => bit_vector(to_signed(32, 16#e9b5dba5#)),   /K_4 => bit_vector(to_signed(32, 16#3956c25b#)),   /K_5 => bit_vector(to_signed(32, 16#59f111f1#)),   /K_6 => bit_vector(to_signed(32, 16#923f82a4#)),   /K_7 => bit_vector(to_signed(32, 16#ab1c5ed5#)),   /K_8 => bit_vector(to_signed(32, 16#d807aa98#)),   /K_9 => bit_vector(to_signed(32, 16#12835b01#)),   0K_10 => bit_vector(to_signed(32, 16#243185be#)),   0K_11 => bit_vector(to_signed(32, 16#550c7dc3#)),   0K_12 => bit_vector(to_signed(32, 16#72be5d74#)),   0K_13 => bit_vector(to_signed(32, 16#80deb1fe#)),   0K_14 => bit_vector(to_signed(32, 16#9bdc06a7#)),   0K_15 => bit_vector(to_signed(32, 16#c19bf174#)),   0K_16 => bit_vector(to_signed(32, 16#e49b69c1#)),   0K_17 => bit_vector(to_signed(32, 16#efbe4786#)),   0K_18 => bit_vector(to_signed(32, 16#0fc19dc6#)),   0K_19 => bit_vector(to_signed(32, 16#240ca1cc#)),   0K_20 => bit_vector(to_signed(32, 16#2de92c6f#)),   0K_21 => bit_vector(to_signed(32, 16#4a7484aa#)),   0K_22 => bit_vector(to_signed(32, 16#5cb0a9dc#)),   0K_23 => bit_vector(to_signed(32, 16#76f988da#)),   0K_24 => bit_vector(to_signed(32, 16#983e5152#)),   0K_25 => bit_vector(to_signed(32, 16#a831c66d#)),   0K_26 => bit_vector(to_signed(32, 16#b00327c8#)),   0K_27 => bit_vector(to_signed(32, 16#bf597fc7#)),   0K_28 => bit_vector(to_signed(32, 16#c6e00bf3#)),   0K_29 => bit_vector(to_signed(32, 16#d5a79147#)),   0K_30 => bit_vector(to_signed(32, 16#06ca6351#)),   0K_31 => bit_vector(to_signed(32, 16#14292967#)),   0K_32 => bit_vector(to_signed(32, 16#27b70a85#)),   0K_33 => bit_vector(to_signed(32, 16#2e1b2138#)),   0K_34 => bit_vector(to_signed(32, 16#4d2c6dfc#)),   0K_35 => bit_vector(to_signed(32, 16#53380d13#)),   0K_36 => bit_vector(to_signed(32, 16#650a7354#)),   0K_37 => bit_vector(to_signed(32, 16#766a0abb#)),   0K_38 => bit_vector(to_signed(32, 16#81c2c92e#)),   0K_39 => bit_vector(to_signed(32, 16#92722c85#)),   0K_40 => bit_vector(to_signed(32, 16#a2bfe8a1#)),   0K_41 => bit_vector(to_signed(32, 16#a81a664b#)),   0K_42 => bit_vector(to_signed(32, 16#c24b8b70#)),   0K_43 => bit_vector(to_signed(32, 16#c76c51a3#)),   0K_44 => bit_vector(to_signed(32, 16#d192e819#)),   0K_45 => bit_vector(to_signed(32, 16#d6990624#)),   0K_46 => bit_vector(to_signed(32, 16#f40e3585#)),   0K_47 => bit_vector(to_signed(32, 16#106aa070#)),   0K_48 => bit_vector(to_signed(32, 16#19a4c116#)),   0K_49 => bit_vector(to_signed(32, 16#1e376c08#)),   0K_50 => bit_vector(to_signed(32, 16#2748774c#)),   0K_51 => bit_vector(to_signed(32, 16#34b0bcb5#)),   0K_52 => bit_vector(to_signed(32, 16#391c0cb3#)),   0K_53 => bit_vector(to_signed(32, 16#4ed8aa4a#)),   0K_54 => bit_vector(to_signed(32, 16#5b9cca4f#)),   0K_55 => bit_vector(to_signed(32, 16#682e6ff3#)),   0K_56 => bit_vector(to_signed(32, 16#748f82ee#)),   0K_57 => bit_vector(to_signed(32, 16#78a5636f#)),   0K_58 => bit_vector(to_signed(32, 16#84c87814#)),   0K_59 => bit_vector(to_signed(32, 16#8cc70208#)),   0K_60 => bit_vector(to_signed(32, 16#90befffa#)),   0K_61 => bit_vector(to_signed(32, 16#a4506ceb#)),   0K_62 => bit_vector(to_signed(32, 16#bef9a3f7#)),   /K_63 => bit_vector(to_signed(32, 16#c67178f2#))   );       type h_vector is record   "    H_0 : bit_vector(31 downto 0);   "    H_1 : bit_vector(31 downto 0);   "    H_2 : bit_vector(31 downto 0);   "    H_3 : bit_vector(31 downto 0);   "    H_4 : bit_vector(31 downto 0);   "    H_5 : bit_vector(31 downto 0);   "    H_6 : bit_vector(31 downto 0);   "    H_7 : bit_vector(31 downto 0);   end record;       constant H : h_vector := (   /H_0 => bit_vector(to_signed(32, 16#6a09e667#)),   /H_1 => bit_vector(to_signed(32, 16#bb67ae85#)),   /H_2 => bit_vector(to_signed(32, 16#3c6ef372#)),   /H_3 => bit_vector(to_signed(32, 16#a54ff53a#)),   /H_4 => bit_vector(to_signed(32, 16#510e527f#)),   /H_5 => bit_vector(to_signed(32, 16#9b05688c#)),   /H_6 => bit_vector(to_signed(32, 16#1f83d9ab#)),   .H_7 => bit_vector(to_signed(32, 16#5be0cd19#))   );5��   .       �       -             b      �      �    -                      �                     �    .                                           �    /                     '                    �    0                     J                    �    1                     m                    �    2                     �                    �    3                     �                    �    4                     �                    �    5                     �                    �    6                                         �    7                     ?                    �    8                     b                    �    9                     �                    �    :                     �                    �    ;                     �                    �    <                     �                    �    =                                         �    >                     9                    �    ?                     ]                    �    @                     �                    �    A                     �                    �    B                     �                    �    C                     �                    �    D                                         �    E                     5                    �    F                     Y                    �    G                     }                    �    H                     �                    �    I                     �                    �    J                     �                    �    K                                         �    L                     1                    �    M                     U                    �    N                     y                    �    O                     �                    �    P                     �                    �    Q                     �                    �    R                     		                    �    S                     -	                    �    T                     Q	                    �    U                     u	                    �    V                     �	                    �    W                     �	                    �    X                     �	                    �    Y                     
                    �    Z                     )
                    �    [                     M
                    �    \                     q
                    �    ]                     �
                    �    ^                     �
                    �    _                     �
                    �    `                                         �    a                     %                    �    b                     I                    �    c                     m                    �    d                     �                    �    e                     �                    �    f                     �                    �    g                     �                    �    h                     !                    �    i                     E                    �    j                     i                    �    k                     �                    �    l                     �                    �    m                     �                    �    n                     �                    �    o                                           �    q                      *                     �    r                      E                     �    s                      u                     �    t                      �                     �    u                      �                     �    v                                           �    w                      5                     �    x                      e                     �    y                      �                     �    z                      �                     �    {                      �                     �    |                      %                     �    }                      V                     �    ~                      �                     �                          �                     �    �                      �                     �    �                                           �    �                      K                     �    �                      |                     �    �                      �                     �    �                      �                     �    �                                           �    �                      @                     �    �                      q                     �    �                      �                     �    �                      �                     �    �                                           �    �                      5                     �    �                      f                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      *                     �    �                      [                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                                           �    �                      P                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                                           �    �                      E                     �    �                      v                     �    �                      �                     �    �                      �                     �    �                      	                     �    �                      :                     �    �                      k                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      /                     �    �                      `                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                      $                     �    �                      U                     �    �                      �                     �    �                      �                     �    �                      �                     �    �                                           �    �                      J                     5�_�               �       ����                                                                                                                                                                                                                                                                                                                ?           8          :                 f�     �   �   �   �          signal clk: bit := '';5��    �                     ."                     5�_�                   �       ����                                                                                                                                                                                                                                                                                                                ?           8          :                 f�     �   �   �   �          signal clk: bit := '0';5��    �                     /"                     5�_�                 4       ����                                                                                                                                                                                                                                                                                                                9                               V       f     �   4   5   �          �   4   6   �           5��    4                      �                     �    4                      �                     �    4                     �                     �    5                                            5�_�               {       ����                                                                                                                                                                                                                                                                                                                7                     	          V       f��     �   z   |   �               K_0 => , 16#428a2f98#)),5��    z                     `                     5�_�                 {       ����                                                                                                                                                                                                                                                                                                                7                     	          V       f��     �   z   |   �              K_0 => ,5��    z                     `                     5�_�                 {       ����                                                                                                                                                                                                                                                                                                                7                     	          V       f��     �   z   |   �              K_0 => "",5��    z                     `                     5�_�                 {       ����                                                                                                                                                                                                                                                                                                                7                     	          V       f��     �   z   |   �              K_0 => ,5��    z                     a                     �    z                     `                     5�_�                 {       ����                                                                                                                                                                                                                                                                                                                7                     	          V       f��     �   z   |   �              K_0 => "",5��    z                     `                     5�_�                 {       ����                                                                                                                                                                                                                                                                                                                7                     	          V       f��     �   z   |   �              K_0 => "00000000",5��    z                     a                     5�_�    	             {       ����                                                                                                                                                                                                                                                                                                                7                     	          V       f��     �   {   |   �    �   z   |   �      "        K_0 => "0000000000000000",5��    z                     i                     5�_�    
          	   {       ����                                                                                                                                                                                                                                                                                                                7                     	          V       f��     �   {   |   �    �   z   |   �      *        K_0 => "000000000000000000000000",5��    z                      q                     5�_�  	              
   {   '    ����                                                                                                                                                                                                                                                                                                                7                     	          V       f��    �   {   |   �    �   z   |   �      2        K_0 => "00000000000000000000000000000000",5��    z   (                  y                     5�_�   �           �   �   n        ����                                                                                                                                                                                                                                                                                                                $           p   !       �   !       V   !    f �
     �   m   o   �      F9a4c116 1e376c08 2748774c 34b0bcb5 391c0cb3 4ed8aa4a 5b9cca4f 682e6ff35��    m                      �                     5�_�   �           �   �          ����                                                                                                                                                                                                                                                                                                                $              	                 v       f �/     �         �      $        if value && (2**i) /= 0 then5��                        �                    5�_�   �           �   �   h   /    ����                                                                                                                                                                                                                                                                                                                           h          o                 f ��     �   g   i   v      6        H_0 => bit_vector(unsigned(16#6a09e667#, 32)),5��    g   /                                        5�_�   q           s   r   k       ����                                                                                                                                                                                                                                                                                                                           d          k                 f ��     �   j   l   r              H_7 => 16#5be0cd19#5��    j                     �                     5�_�   g   i       k   h   d       ����                                                                                                                                                                                                                                                                                                                           k          d          V       f �9     �   c   e   r      V        H_0 => 6a09e667bb67ae85 3c6ef372 a54ff53a 510e527f 9b05688c 1f83d9ab 5be0cd19,5��    c                     �                     5�_�   h   j           i   d       ����                                                                                                                                                                                                                                                                                                                           k          d          V       f �;     �   c   e   r              H_0 => 6a09e667,5��    c          >           �      >               5�_�   i               j   f       ����                                                                                                                                                                                                                                                                                                                           k          d          V       f �A     �   e   g   r             ,5��    e                     �                     5�_�   Z           \   [   b        ����                                                                                                                                                                                                                                                                                                                                      a           V        f �     �   b   c   h    �   b   c   h   8           H_8 : integer;           H_9 : integer;           H_10 : integer;           H_11 : integer;           H_12 : integer;           H_13 : integer;           H_14 : integer;           H_15 : integer;           H_16 : integer;           H_17 : integer;           H_18 : integer;           H_19 : integer;           H_20 : integer;           H_21 : integer;           H_22 : integer;           H_23 : integer;           H_24 : integer;           H_25 : integer;           H_26 : integer;           H_27 : integer;           H_28 : integer;           H_29 : integer;           H_30 : integer;           H_31 : integer;           H_32 : integer;           H_33 : integer;           H_34 : integer;           H_35 : integer;           H_36 : integer;           H_37 : integer;           H_38 : integer;           H_39 : integer;           H_40 : integer;           H_41 : integer;           H_42 : integer;           H_43 : integer;           H_44 : integer;           H_45 : integer;           H_46 : integer;           H_47 : integer;           H_48 : integer;           H_49 : integer;           H_50 : integer;           H_51 : integer;           H_52 : integer;           H_53 : integer;           H_54 : integer;           H_55 : integer;           H_56 : integer;           H_57 : integer;           H_58 : integer;           H_59 : integer;           H_60 : integer;           H_61 : integer;           H_62 : integer;           H_63 : integer;5��    b               8       �              >      5�_�   V       W   Y   X           ����                                                                                                                                                                                                                                                                                                                           _   	                 V   	    f ��     �         g      *    type k_vector is record K_0 : integer;5��                             	              5�_�   V           X   W           ����                                                                                                                                                                                                                                                                                                                           `   	          	       V   	    f ��     �         g              K_0 : bit_vector;�                        K_1 : bit_vector;�                        K_2 : bit_vector;�                        K_3 : bit_vector;�                        K_4 : bit_vector;�                        K_5 : bit_vector;�                        K_6 : bit_vector;�                        K_7 : bit_vector;�                        K_8 : bit_vector;�                         K_9 : bit_vector;�      !                  K_10 : bit_vector;�       "                  K_11 : bit_vector;�   !   #                  K_12 : bit_vector;�   "   $                  K_13 : bit_vector;�   #   %                  K_14 : bit_vector;�   $   &                  K_15 : bit_vector;�   %   '                  K_16 : bit_vector;�   &   (                  K_17 : bit_vector;�   '   )                  K_18 : bit_vector;�   (   *                  K_19 : bit_vector;�   )   +                  K_20 : bit_vector;�   *   ,                  K_21 : bit_vector;�   +   -                  K_22 : bit_vector;�   ,   .                  K_23 : bit_vector;�   -   /                  K_24 : bit_vector;�   .   0                  K_25 : bit_vector;�   /   1                  K_26 : bit_vector;�   0   2                  K_27 : bit_vector;�   1   3                  K_28 : bit_vector;�   2   4                  K_29 : bit_vector;�   3   5                  K_30 : bit_vector;�   4   6                  K_31 : bit_vector;�   5   7                  K_32 : bit_vector;�   6   8                  K_33 : bit_vector;�   7   9                  K_34 : bit_vector;�   8   :                  K_35 : bit_vector;�   9   ;                  K_36 : bit_vector;�   :   <                  K_37 : bit_vector;�   ;   =                  K_38 : bit_vector;�   <   >                  K_39 : bit_vector;�   =   ?                  K_40 : bit_vector;�   >   @                  K_41 : bit_vector;�   ?   A                  K_42 : bit_vector;�   @   B                  K_43 : bit_vector;�   A   C                  K_44 : bit_vector;�   B   D                  K_45 : bit_vector;�   C   E                  K_46 : bit_vector;�   D   F                  K_47 : bit_vector;�   E   G                  K_48 : bit_vector;�   F   H                  K_49 : bit_vector;�   G   I                  K_50 : bit_vector;�   H   J                  K_51 : bit_vector;�   I   K                  K_52 : bit_vector;�   J   L                  K_53 : bit_vector;�   K   M                  K_54 : bit_vector;�   L   N                  K_55 : bit_vector;�   M   O                  K_56 : bit_vector;�   N   P                  K_57 : bit_vector;�   O   Q                  K_58 : bit_vector;�   P   R                  K_59 : bit_vector;�   Q   S                  K_60 : bit_vector;�   R   T                  K_61 : bit_vector;�   S   U                  K_62 : bit_vector;�   T   V                  K_63 : bit_vector;�   X   Z                  H_0 : bit_vector;�   Y   [                  H_1 : bit_vector;�   Z   \                  H_2 : bit_vector;�   [   ]                  H_3 : bit_vector;�   \   ^                  H_4 : bit_vector;�   ]   _                  H_5 : bit_vector;�   ^   `                  H_6 : bit_vector;�   _   a                  H_7 : bit_vector;5��                     
   *             
       �                     
   D             
       �                     
   ^             
       �                     
   x             
       �                     
   �             
       �                     
   �             
       �                     
   �             
       �                     
   �             
       �                     
   �             
       �                     
                
       �                     
   /             
       �                      
   J             
       �    !                 
   e             
       �    "                 
   �             
       �    #                 
   �             
       �    $                 
   �             
       �    %                 
   �             
       �    &                 
   �             
       �    '                 
                
       �    (                 
   "             
       �    )                 
   =             
       �    *                 
   X             
       �    +                 
   s             
       �    ,                 
   �             
       �    -                 
   �             
       �    .                 
   �             
       �    /                 
   �             
       �    0                 
   �             
       �    1                 
                
       �    2                 
   0             
       �    3                 
   K             
       �    4                 
   f             
       �    5                 
   �             
       �    6                 
   �             
       �    7                 
   �             
       �    8                 
   �             
       �    9                 
   �             
       �    :                 
                
       �    ;                 
   #             
       �    <                 
   >             
       �    =                 
   Y             
       �    >                 
   t             
       �    ?                 
   �             
       �    @                 
   �             
       �    A                 
   �             
       �    B                 
   �             
       �    C                 
   �             
       �    D                 
                
       �    E                 
   1             
       �    F                 
   L             
       �    G                 
   g             
       �    H                 
   �             
       �    I                 
   �             
       �    J                 
   �             
       �    K                 
   �             
       �    L                 
   �             
       �    M                 
   	             
       �    N                 
   $             
       �    O                 
   ?             
       �    P                 
   Z             
       �    Q                 
   u             
       �    R                 
   �             
       �    S                 
   �             
       �    T                 
   �             
       �    X                 
   	             
       �    Y                 
   +	             
       �    Z                 
   E	             
       �    [                 
   _	             
       �    \                 
   y	             
       �    ]                 
   �	             
       �    ^                 
   �	             
       �    _                 
   �	             
       5�_�   L           N   M      
    ����                                                                                                                                                                                                                                                                                                                              
          
          
    f �9     �          ]   	           H_1 : integer;           H_2 : integer;           H_3 : integer;           H_4 : integer;           H_5 : integer;           H_6 : integer;           H_7 : integer;           H_8 : integer;           H_9 : integer;5��       
                 =                    �       
                 T                    �       
                 k                    �       
                 �                    �       
                 �                    �       
                 �                    �       
                 �                    �       
                 �                    �       
                 �                    5�_�   J           L   K          ����                                                                                                                                                                                                                                                                                                                                                      f ��     �             �                       H_0 : integer;5��                          3                     5�_�   /           1   0      !    ����                                                                                                                                                                                                                                                                                                                                                             f �\     �               -        haso : out bit_vector(255downto 0 ) ;5��       !                  �                      5�_�                          ����                                                                                                                                                                                                                                                                                                                                                             f �K     �               1        msgi : in bit_vect  r (5 1 1 downto 0 ) ;5��                         V                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f �K     �               0        msgi : in bit_vect   (5 1 1 downto 0 ) ;5��                         W                      5��