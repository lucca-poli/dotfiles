Vim�UnDo� ng^���"����/D��o75	�q�
t/   Z           wait for CLOCK_PERIOD;   I         �       �   �   �    fǺ    _�                     	        ����                                                                                                                                                                                                                                                                                                                            	                      V        f��     �         M    �   	   
   M    �      	          C            clk : in bit;                            -- Clock input   A            rst : in bit;                          -- Reset input   F            count : out integer       -- 6-bit count output (64 steps)5��                          �       �               �                          �               �       5�_�                    	       ����                                                                                                                                                                                                                                                                                                                            	                           f��     �   	      P              done: out bit;   B        count : out natural       -- 6-bit count output (64 steps)�      
   P      J        clk, rst, start: in bit;                            -- Clock input5��                         �                      �    	                     �                      �    
                     	                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         P      -    signal rst : bit := '0';  -- Reset signal5��                        �                    �                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         P      -    signal clk : bit := '0';  -- Clock signal5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         P      /    signal clk,  : bit := '0';  -- Clock signal�         P    5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         P      2    signal clk, rst : bit := '0';  -- Clock signal5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f�     �         P      8    signal clk, rst, done : bit := '0';  -- Clock signal5��                         �                     5�_�      	                     ����                                                                                                                                                                                                                                                                                                                            	                           f�     �                *    signal  : bit := '0';  -- Reset signal5��                          �      +               5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                            	                           f�     �         O          component counter_6bit5��                        �                     5�_�   	              
   !   	    ����                                                                                                                                                                                                                                                                                                                            !   	       !          v       f�!     �       "   O          dut: counter_6bit�   !   "   O    5��        	                 H                    5�_�   
                 $        ����                                                                                                                                                                                                                                                                                                                            !   	       !          v       f�*     �   "   $   M                  clk => clk,�   #   $                      rst => rst,               count => count5��    #                      �      3               �    "                     w                     �    "                     k                    �    "                     l                     �    "                      k                     5�_�                    $       ����                                                                                                                                                                                                                                                                                                                            !   	       !          v       f�,     �   !   #   K              port map (clk, rst);�   !   #   L              port map (   );�   "   $   M          );�   #   %   M      
        );5��    #                     m                     �    #                      l                     �    "                      k                     �    !                     j                     �    !                     j                     �    !                     p                     �    !                    o                    �    !                    o                    �    !                    o                    �    !                    t                    �    !                     u                     �    !                    t                    �    !                    t                    �    !                 	   t             	       �    !   $                  |                     �    !   #                 {                    �    !   #                 {                    �    !   #              	   {             	       �    !   +                  �                     �    !   *                  �                     �    !   )                 �                    �    !   )                 �                    �    !   )                 �                    5�_�                    E       ����                                                                                                                                                                                                                                                                                                                            !   	       !          v       f�X     �   E   H   L              �   E   G   K    5��    E                                    	       �    E                                           �    E                                   	       �    F                                           5�_�                    G        ����                                                                                                                                                                                                                                                                                                                            !   	       !          v       f�Y     �   G   I   M    �   G   H   M    5��    G                                           5�_�                    G        ����                                                                                                                                                                                                                                                                                                                            !   	       !          v       f�Z     �   F   G           5��    F                                           5�_�                           ����                                                                                                                                                                                                                                                                                                                            !   	       !          v       f�p     �         M    �         M    5��                          �              @       5�_�                           ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       f�s     �         N      ?    signal clk, rst, start, done : bit := '0';  -- Clock signal5��              
                 
               5�_�                           ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       f�v     �         N      5    signal start, done : bit := '0';  -- Clock signal5��                                              5�_�                           ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       f�y     �         N      .    signal start: bit := '0';  -- Clock signal5��                                            5�_�                           ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       f�|     �         N      ?    signal clk, rst, start, done : bit := '0';  -- Clock signal5��                         �                     5�_�                    1       ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       fҌ     �   0   2   O              �   0   2   N    5��    0                      �              	       �    0                     �                     �    0   
                  �                     �    0   	                  �                     �    0                    �                    �    0                    �                    �    0                 	   �             	       5�_�                    1       ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       fґ     �   0   2   O              start <= 5��    0                     �                     5�_�                    1       ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       fґ     �   0   2   O              start <= ''5��    0                                           5�_�                    1       ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       fғ     �   0   2   O              start <= '0'5��    0                                          5�_�                    #       ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       fҡ     �   "   $   O    �   #   $   O    5��    "                      �              1       5�_�                    #       ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       fҢ     �   "   $   P      0        port map (clk, rst, start, done, count);5��    "                    �                    5�_�                    #       ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       fҩ     �   "   $   P      3        generic map (clk, rst, start, done, count);5��    "                    �                    �    "                    �                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            "   	       "          v       f��     �         P    �         P    5��                          �               /       5�_�                           ����                                                                                                                                                                                                                                                                                                                                      
                 f��     �         S              MAX_COUNT: natural       );�      	   S          generic(5��                         �                      �                         �                      �    	                     �                      5�_�                    &       ����                                                                                                                                                                                                                                                                                                                                      
                 f��     �   %   '   S              generic map (8);5��    %                     �                     5�_�                     1   E    ����                                                                                                                                                                                                                                                                                                                                      
                 f��     �   0   2   S      V        "Did not proceed to 1, count is " & integer'image(to_integer(unsigned(count)))5��    0   E                  �                     5�_�      !               1   E    ����                                                                                                                                                                                                                                                                                                                                      
                 f��     �   0   2   S      N        "Did not proceed to 1, count is " & integer'image(to_integer((count)))5��    0   E                  �                     5�_�       "           !   1   J    ����                                                                                                                                                                                                                                                                                                                                      
                 f��     �   0   2   S      M        "Did not proceed to 1, count is " & integer'image(to_integer(count)))5��    0   J                  �                     5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                                      
                 f��     �         S      .    signal count : integer;  -- Input stimulus5��                        l                    �                         q                     �                         p                     �                         o                     �                         n                     �                         m                     �                        l                    �                        l                    �                        l                    5�_�   "   $           #   1   :    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   0   2   S      L        "Did not proceed to 1, count is " & integer'image(to_integer(count))5��    0   :       
           �      
               5�_�   #   %           $   1   :    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   0   2   S      B        "Did not proceed to 1, count is " & integer'image((count))5��    0   :                  �                     5�_�   $   &           %   1   ?    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   0   2   S      A        "Did not proceed to 1, count is " & integer'image(count))5��    0   ?                  �                     5�_�   %   '           &   7   :    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   6   8   S      V        "Did not proceed to 2, count is " & integer'image(to_integer(unsigned(count)))5��    6   :                  �                     5�_�   &   (           '   7   9    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   6   8   S      C        "Did not proceed to 2, count is " & integer'image((count)))5��    6   9                  �                     5�_�   '   )           (   7   ?    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   6   8   S      B        "Did not proceed to 2, count is " & integer'image(count)))5��    6   ?                  �                     5�_�   (   *           )   7   ?    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   6   8   S      A        "Did not proceed to 2, count is " & integer'image(count))5��    6   ?                  �                     5�_�   )   +           *   <   :    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   ;   =   S      V        "Did not proceed to 3, count is " & integer'image(to_integer(unsigned(count)))5��    ;   :                  6                     5�_�   *   ,           +   <   :    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   ;   =   S      C        "Did not proceed to 3, count is " & integer'image((count)))5��    ;   :                  6                     5�_�   +   -           ,   <   ?    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   ;   =   S      B        "Did not proceed to 3, count is " & integer'image(count)))5��    ;   ?                  ;                     5�_�   ,   .           -   <   ?    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   ;   =   S      A        "Did not proceed to 3, count is " & integer'image(count))5��    ;   ?                  ;                     5�_�   -   /           .   A   :    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   @   B   S      W        "Did not proceed to 4, count is " & integer'image(to_integer(unsigned(count))) 5��    @   :                  �                     5�_�   .   0           /   A   ?    ����                                                                                                                                                                                                                                                                                                                                      
                 f�     �   @   B   S      C        "Did not proceed to 4, count is " & integer'image(count))) 5��    @   ?                  �                     5�_�   /   1           0   A   ?    ����                                                                                                                                                                                                                                                                                                                                      
                 f�    �   @   B   S      B        "Did not proceed to 4, count is " & integer'image(count)) 5��    @   ?                  �                     5�_�   0   2           1           ����                                                                                                                                                                                                                                                                                                                            K   ?       F   $       V   ?    f�D     �               S   library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity counter_tb is end;       (architecture Behavioral of counter_tb is       component counter_generic           generic(               MAX_COUNT: natural   
        );           port (   N            clk, rst, start: in bit;                            -- Clock input               done: out bit;   F            count : out natural       -- 6-bit count output (64 steps)   
        );       end component;       J    constant CLOCK_PERIOD : time := 20 ns;  -- Clock period (e.g., 50 MHz)       8    signal clk, rst, done : bit := '0';  -- Clock signal   .    signal start: bit := '1';  -- Clock signal   .    signal count : natural;  -- Input stimulus       begin       -- Clock process       clk_process: process   	    begin           clk <= '0';   "        wait for CLOCK_PERIOD / 2;           while true loop               clk <= not clk;   &            wait for CLOCK_PERIOD / 2;           end loop;       end process clk_process;           -- DUT instantiation       dut: counter_generic           generic map (8)   0        port map (clk, rst, start, done, count);           -- Stimulus process       stim: process   	    begin       6        assert false report "BOT count" severity note;               wait for CLOCK_PERIOD;            assert count = 1 report    @        "Did not proceed to 1, count is " & integer'image(count)           severity error;               wait for CLOCK_PERIOD;           start <= '0';            assert count = 2 report    @        "Did not proceed to 2, count is " & integer'image(count)           severity error;               wait for CLOCK_PERIOD;            assert count = 3 report    @        "Did not proceed to 3, count is " & integer'image(count)           severity error;               wait for CLOCK_PERIOD;            assert count = 4 report    A        "Did not proceed to 4, count is " & integer'image(count)            severity error;               wait for CLOCK_PERIOD;       $        rst <= '1';  -- Assert reset   7        wait for CLOCK_PERIOD;  -- Hold reset for 20 ns   ?        assert count = 0 report "Did not reset" severity error;   &        rst <= '0';  -- Deassert reset   7        wait for CLOCK_PERIOD;  -- Hold reset for 20 ns   A        assert count = 1 report "Did not proceed" severity error;               wait for CLOCK_PERIOD;       6        assert false report "EOT count" severity note;               wait;       end process stim;   end Behavioral;5�5�_�   1   3           2   1   ,    ����                                                                                                                                                                                                                                                                                                                            K   ?       F   $       V   ?    f��     �   0   2   S      @        "Did not proceed to 1, count is " & integer'image(count)5��    0   ,                  �                     5�_�   2   4           3   1   ,    ����                                                                                                                                                                                                                                                                                                                            K   ?       F   $       V   ?    f��     �   0   2   S      ,        "Did not proceed to 1, count is " & 5��    0   ,                  �                     �    0   -                  �                     �    0   ,                  �                     �    0   +                 �                    �    0   -                 �                    5�_�   3   5           4   1   -    ����                                                                                                                                                                                                                                                                                                                            K   ?       F   $       V   ?    f��     �   1   3   S    5��    1                      �              	       �    1                      �                     5�_�   4   6           5   2        ����                                                                                                                                                                                                                                                                                                                            L   ?       G   $       V   ?    f��     �   1   3   T       �   2   3   T    5��    1                      �                     5�_�   5   7           6   2        ����                                                                                                                                                                                                                                                                                                                            L   ?       G   $       V   ?    f��     �   1   3   T      integer'image(count)5��    1                      �                     5�_�   6   8           7   2       ����                                                                                                                                                                                                                                                                                                                            L   ?       G   $       V   ?    f��     �   1   3   T              integer'image(count)5��    1                     �                     �    1   	                 �                    5�_�   7   9           8   2       ����                                                                                                                                                                                                                                                                                                                            L   ?       G   $       V   ?    f��     �   1   3   T      *        "count is: " &integer'image(count)5��    1                     �                     5�_�   8   :           9   1       ����                                                                                                                                                                                                                                                                                                                            L   ?       G   $       V   ?    f��     �   0   2   T      .        "Did not proceed to 1, count is " &LF&5��    0                     �                     5�_�   9   ;           :   2   +    ����                                                                                                                                                                                                                                                                                                                            L   ?       G   $       V   ?    f��     �   1   4   T      +        "count is: " & integer'image(count)5��    1   +                                       �    1   ,                                     �    1   0                               	       5�_�   :   <           ;   3       ����                                                                                                                                                                                                                                                                                                                            M   ?       H   $       V   ?    f��     �   2   4   U              5��    2                                          5�_�   ;   =           <   3   	    ����                                                                                                                                                                                                                                                                                                                            M   ?       H   $       V   ?    f��     �   2   4   U      
        ""5��    2   	               
                 
       5�_�   <   >           =   3       ����                                                                                                                                                                                                                                                                                                                            M   ?       H   $       V   ?    f��     �   2   4   U              "start is: "5��    2                                          �    2                                          �    2                 	                	       �    2                     &                     �    2                     %                     �    2                     $                     �    2                     #                     �    2                    "                    �    2                    "                    �    2                    "                    5�_�   =   ?           >   3        ����                                                                                                                                                                                                                                                                                                                            M   ?       H   $       V   ?    f�     �   2   4   U               "start is: " & bit'image5��    2                      '                     5�_�   >   @           ?   3   !    ����                                                                                                                                                                                                                                                                                                                            M   ?       H   $       V   ?    f�     �   2   4   U      "        "start is: " & bit'image()5��    2   !                  (                     �    2   #                  *                     �    2   "                  )                     �    2   !                 (                    �    2   !                 (                    �    2   !                 (                    5�_�   ?   A           @   9   %    ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    f�     �   9   <   U    �   9   :   U    5��    9                      �              Y       5�_�   @   B           A   @       ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    f�!     �   @   C   W    �   @   A   W    5��    @                      �              Y       5�_�   A   D           B   G       ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    f�"     �   G   J   Y    �   G   H   Y    5��    G                      �              Y       5�_�   B   E   C       D   9       ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    f�@     �   8   :   [      @        "Did not proceed to 2, count is " & integer'image(count)5��    8                     �                     5�_�   D   F           E   9       ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    f�E     �   8   :   [      5        "Did not proceed to 2" & integer'image(count)5��    8                    �                    5�_�   E   G           F   @       ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    f�Q     �   ?   A   [      @        "Did not proceed to 3, count is " & integer'image(count)5��    ?                     �                     �    ?                    �                    5�_�   F   H           G   G       ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    f�T    �   F   H   [      A        "Did not proceed to 4, count is " & integer'image(count) 5��    F                     g                     �    F                    h                    5�_�   G   I           H   3        ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    fղ     �   3   5   [    5��    3                      /              	       5�_�   H   J           I   4       ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    fճ     �   3   5   \              5��    3                     7                     5�_�   I   K           J   4   	    ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    fմ     �   3   5   \      
        ""5��    3   	                  8                     5�_�   J   L           K   4       ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    fչ     �   3   5   \              "rst is: "5��    3                     A                     5�_�   K   M           L   4       ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    fտ     �   3   5   \              "rst is: " & bit'image5��    3                     M                     5�_�   L   N           M   4       ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    fտ     �   3   5   \               "rst is: " & bit'image()5��    3                     N                     �    3                    N                    5�_�   M   O           N   4   #    ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    f��     �   3   5   \      #        "rst is: " & bit'image(rst)5��    3   #                  R                     �    3   #                  R                     5�_�   N   P           O   3   '    ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    f��    �   2   4   \      '        "start is: " & bit'image(start)5��    2   '                  .                     5�_�   O   Q           P          ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    f��    �         \      .    signal count : natural;  -- Input stimulus5��                         s                     �                        t                    5�_�   P   R           Q          ����                                                                                                                                                                                                                                                                                                                                                             f�D     �         \      3    signal count : natural := 0;  -- Input stimulus5��                         s                     5�_�   Q   S           R          ����                                                                                                                                                                                                                                                                                                                                                             f�K     �         \      8    signal clk, rst, done : bit := '0';  -- Clock signal5��                                              5�_�   R   T           S          ����                                                                                                                                                                                                                                                                                                                                                             f�K     �         \      6    signal clk, rstdone : bit := '0';  -- Clock signal5��                                              5�_�   S   U           T          ����                                                                                                                                                                                                                                                                                                                                                             f�O     �         \    �         \    5��                          R              /       5�_�   T   V           U          ����                                                                                                                                                                                                                                                                                                                                                             f�P     �         ]      .    signal start: bit := '1';  -- Clock signal5��                        ]                    5�_�   U   W           V          ����                                                                                                                                                                                                                                                                                                                                                             f�U    �         ]      -    signal done: bit := '1';  -- Clock signal5��                         f                     5�_�   V   X           W   0       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   0   2   ^              �   0   2   ]    5��    0                      �              	       �    0                     �                     �    0   
                  �                     �    0   	                  �                     �    0                    �                    �    0                    �                    �    0                 
   �             
       �    0                     �                     5�_�   W   Y           X   1       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   0   2   ^              start <= 5��    0                     �                     5�_�   X   Z           Y   1       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   0   2   ^              start <= ''5��    0                     �                     5�_�   Y   [           Z   1       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   0   2   ^              start <= '1;'5��    0                     �                     5�_�   Z   \           [   1       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   0   2   ^              start <= '1'�   1   2   ^    5��    0                     �                     5�_�   [   ]           \   1       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   1   3   ^    �   1   2   ^    5��    1                      �                     5�_�   \   ^           ]   2       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   1   3   _              start <= '1';5��    1                    �                    �    1                     �                     5�_�   ]   _           ^   2       ����                                                                                                                                                                                                                                                                                                                                                             f��    �   1   2                   <= '1';5��    1                      �                     5�_�   ^   `           _   #        ����                                                                                                                                                                                                                                                                                                                                       ^           V        f��     �   #   %   ^    �   #   $   ^    5��    #                      �                     5�_�   _   a           `          ����                                                                                                                                                                                                                                                                                                                            #                    V       f�     �             
       -- Clock process       clk_process: process   	    begin           clk <= '0';   "        wait for CLOCK_PERIOD / 2;           while true loop               clk <= not clk;   &            wait for CLOCK_PERIOD / 2;           end loop;       end process clk_process;5��           
               �      �               5�_�   `   b           a          ����                                                                                                                                                                                                                                                                                                                                                V       f�     �         U          clk <= not clk after 5 ns;5��                        �                    �                         �                     �                        �                    �                        �                    �                        �                    5�_�   a   c           b   T       ����                                                                                                                                                                                                                                                                                                                                                V       f�?     �   S   U   U          end process stim;5��    S                     B	                     5�_�   b   d           c   T       ����                                                                                                                                                                                                                                                                                                                                                V       f�@     �   S   U   U          end process ;5��    S                     A	                     5�_�   c   e           d   "       ����                                                                                                                                                                                                                                                                                                                                                V       f�E    �   !   #   U          stim: process5��    !                     o                     5�_�   d   f           e           ����                                                                                                                                                                                                                                                                                                                                                V       f�     �         T    �         T    �                &    clk <= not clk after CLOCK_PERIOD;5��                          �      '               �                          �              H       5�_�   e   g           f          ����                                                                                                                                                                                                                                                                                                                                          F       V       f�     �         U      G    clock <= not clock after half_period when finished /= '1' else '0';5��                        �                    5�_�   f   h           g          ����                                                                                                                                                                                                                                                                                                                                          F       V       f�
     �         U      E    clk <= not clock after half_period when finished /= '1' else '0';5��                        �                    5�_�   g   i           h          ����                                                                                                                                                                                                                                                                                                                                          F       V       f�     �         U      C    clk <= not clk after half_period when finished /= '1' else '0';5��                         �                     5�_�   h   j           i          ����                                                                                                                                                                                                                                                                                                                                          F       V       f�     �         U      8    clk <= not clk after  when finished /= '1' else '0';5��                         �                     5�_�   i   k           j          ����                                                                                                                                                                                                                                                                                                                                          F       V       f�     �         U      :    clk <= not clk after () when finished /= '1' else '0';5��                         �                     �                        �                    �                        �                    �                        �                    �                        �                    �                        �                    5�_�   j   l           k      )    ����                                                                                                                                                                                                                                                                                                                                          F       V       f�     �         W      
    signal�         V          �         U    5��                          �                     �                          �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    �                         �                     �                         �                     �                         �                     �                        �                    �                        �                    �                     	   �             	       �                     	   �             	       5�_�   k   m           l          ����                                                                                                                                                                                                                                                                                                                                          F       V       f�      �         W          signal finished: bit := 5��                         �                     5�_�   l   n           m          ����                                                                                                                                                                                                                                                                                                                                          F       V       f�      �         W          signal finished: bit := ''5��                         �                     5�_�   m   p           n          ����                                                                                                                                                                                                                                                                                                                                          F       V       f�!     �         W          signal finished: bit := '0'5��                         �                     5�_�   n   q   o       p   P        ����                                                                                                                                                                                                                                                                                                                                          F       V       f�1     �   P   R   X              �   P   R   W    5��    P                      	                     �    P                      	                     5�_�   p   r           q   Q   
    ����                                                                                                                                                                                                                                                                                                                                          F       V       f�4     �   P   Q                  fin5��    P                      	                     5�_�   q   s           r   Q   
    ����                                                                                                                                                                                                                                                                                                                                          F       V       f�5     �   Q   S   X              �   Q   S   W    5��    Q                      +	              	       �    Q                     3	                     �    Q   
                  5	                     �    Q   	                  4	                     �    Q                    3	                    �    Q                    3	                    �    Q                    3	                    5�_�   r   t           s   R       ����                                                                                                                                                                                                                                                                                                                                          F       V       f�9     �   Q   S   X              finished <= 5��    Q                     ?	                     5�_�   s   u           t   R       ����                                                                                                                                                                                                                                                                                                                                          F       V       f�9     �   Q   S   X              finished <= ''5��    Q                     @	                     5�_�   t   v           u   R       ����                                                                                                                                                                                                                                                                                                                                          F       V       f�;   	 �   Q   S   X              finished <= '1'5��    Q                     B	                     5�_�   u   w           v      	    ����                                                                                                                                                                                                                                                                                                                               	                 v       f'�   
 �          X          dut: counter_generic�          X    5��       	                 ?                    5�_�   v   x           w   
   
    ����                                                                                                                                                                                                                                                                                                                                      X          V       f@;     �   	      X      
        );5��    	   	                  �                      5�_�   w   y           x   
   	    ����                                                                                                                                                                                                                                                                                                                                      X          V       f@D    �   	      X      	        )5��    	   	                  �                      5�_�   x   z           y   *       ����                                                                                                                                                                                                                                                                                                                                      X          V       fB�     �   )   *                  start <= '1';5��    )                                           5�_�   y   {           z   2       ����                                                                                                                                                                                                                                                                                                                                      W          V       fB�     �   1   3   W              start <= '0';5��    1                    0                    5�_�   z   |           {   *       ����                                                                                                                                                                                                                                                                                                                                      W          V       fB�     �   )   +   W    �   *   +   W    5��    )                                           5�_�   {   ~           |   *       ����                                                                                                                                                                                                                                                                                                                                      X          V       fB�    �   )   +   X              start <= '1';5��    )                    1                    5�_�   |      }       ~   ;       ����                                                                                                                                                                                                                                                                                                                                      X          V       fB�    �   :   <   X    �   ;   <   X    5��    :                                            5�_�   ~   �              K       ����                                                                                                                                                                                                                                                                                                                                      Y          V       fB�     �   K   M   Y    �   K   L   Y    5��    K                                           5�_�      �           �   L       ����                                                                                                                                                                                                                                                                                                                                      Z          V       fB�    �   K   M   Z              start <= '0';5��    K                                        5�_�   �   �           �   I        ����                                                                                                                                                                                                                                                                                                                                                             fǰ     �   I   K   Z    �   I   J   Z    5��    I                      �                     5�_�   �   �           �   J       ����                                                                                                                                                                                                                                                                                                                                                             fǰ     �   J   L   [    �   J   K   [    5��    J                                           5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                                                             fǰ     �   K   M   \    �   K   L   \    5��    K                                            5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                                                             fǰ     �   L   N   ]    �   L   M   ]    5��    L                      ?                     5�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                                                             fǰ     �   M   O   ^    �   M   N   ^    5��    M                      ^                     5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                                                             fǱ     �   N   P   _    �   N   O   _    5��    N                      }                     5�_�   �   �           �   O       ����                                                                                                                                                                                                                                                                                                                                                             fǱ     �   O   Q   `    �   O   P   `    5��    O                      �                     5�_�   �   �           �   P       ����                                                                                                                                                                                                                                                                                                                                                             fǳ     �   O   P                  wait for CLOCK_PERIOD;5��    O                      �                     5�_�   �   �           �   K        ����                                                                                                                                                                                                                                                                                                                                                             fǶ     �   J   K                  wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;5��    J                            �               5�_�   �   �           �   J        ����                                                                                                                                                                                                                                                                                                                                                             fǷ     �   I   J                  wait for CLOCK_PERIOD;5��    I                      �                     5�_�   �               �   I       ����                                                                                                                                                                                                                                                                                                                                                             fǹ    �   H   J   Z              wait for CLOCK_PERIOD;5��    H                     �                     5�_�   |           ~   }   B       ����                                                                                                                                                                                                                                                                                                                                      X          V       fB�    �   A   C   X               assert count = 7 report 5��    A                                        5�_�   n           p   o   Q       ����                                                                                                                                                                                                                                                                                                                                          F       V       f�/     �   Q   R   W       5��    Q                      +	              	       �    Q                      +	                     5�_�   B           D   C   9       ����                                                                                                                                                                                                                                                                                                                            3   %       2   %       V   %    f�3     �   8   :   [      5        "Did not proceed to 2" & integer'image(count)5��    8                     �                     5��