Vim�UnDo� *} �d��IՔ���X�;5t~l�fK�6����   f   entity interface_hcsr04_uc is                               fs    _�                              ����                                                                                                                                                                                                                                                                                                                                                             fs    �                /architecture fsm_arch of interface_hcsr04_uc is�                end interface_hcsr04_uc;�         f      entity interface_hcsr04_uc is 5��                        3                     �                        �                    �                        
                    5��