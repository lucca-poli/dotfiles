Vim�UnDo� ���'CV�M�.Ϭ������%(~(*�AjI   �   +    r(31) <= A(31) xor B(31) xor carry(31);   �         1       1   1   1    f��    _�                             ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�'     �         '    5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�*     �         (    5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�+     �         )       �        )    5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�-     �                 antonio.seabra@usp.br5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�H     �         )       �        )    5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�I     �                 antonio.seabra@usp.br5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�P     �         )       �        )    5��                                           #      5�_�      	                      ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�Q     �                 5��                          #                     5�_�                 	           ����                                                                                                                                                                                                                                                                                                                                                 V       f�i    �                 library IEEE;   "use IEEE.NUMERIC_BIT_UNSIGNED.ALL;       entity sigma0 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end sigma0;       architecture arch5 of sigma0 is   begin   0    q <= (x ror 7) xor (x ror 18) xor (x srl 3);   
end arch5;       library IEEE;   "use IEEE.NUMERIC_BIT_UNSIGNED.ALL;       entity sigma1 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end sigma1;       architecture arch6 of sigma1 is   begin   2    q <= (x ror 17) xor (x ror 19) xor (x srl 10);   
end arch6;    5��                                   $              5�_�   	                        ����                                                                                                                                                                                                                                                                                                                            �   G       �   G       V   G    f6�    �  &  (          end somadorarch;�   �   �          &architecture somadorarch of somador is�   �   �          end somador;�   �   �          entity somador is�   �   �          	--somador�   �   �          ^        inst13: somador port map (a => hout, b => x"5be0cd19",  soma => haso(255 downto 224));�   �   �          ^        inst12: somador port map (a => gout, b => x"1f83d9ab",  soma => haso(223 downto 192));�   �   �          ^        inst11: somador port map (a => fout, b => x"9b05688c",  soma => haso(191 downto 160));�   �   �          ^        inst10: somador port map (a => eout, b => x"510e527f",  soma => haso(159 downto 128));�   �   �          \        inst9: somador port map (a => dout, b => x"a54ff53a",  soma => haso(127 downto 96));�   �   �          [        inst8: somador port map (a => cout, b => x"3c6ef372",  soma => haso(95 downto 64));�   �   �          [        inst7: somador port map (a => bout, b => x"bb67ae85",  soma => haso(63 downto 32));�   �   �          Z        inst6: somador port map (a => aout, b => x"6a09e667",  soma => haso(31 downto 0));�   �   �          E        	sum: somador port map(a => waux, b => kaux, soma => kpwaux);�   �   �          2        	inst5: somador port map(y4, W(i-16), y5);�   �   �          -        	inst4: somador port map(y3, y2, y4);�   �   �          1        	inst3: somador port map(y1, W(i-7), y3);�        '      component somador is5��       
              
   �             
       �    �                 
   �             
       �    �                 
   �             
       �    �                 
                
       �    �                 
                
       �    �                 
   �             
       �    �                 
                
       �    �                 
   x             
       �    �                 
   �             
       �    �                 
   8             
       �    �                 
   �             
       �    �                 
   �             
       �    �                 
   ^             
       �    �                 
   �             
       �    �                 
   �             
       �    �                 
   N             
       �    �                 
   h             
       �    �                 
   z             
       �    &                
   �'             
       5�_�                            ����                                                                                                                                                                                                                                                                                                                            �   G       �   G       V   G    f6�    �                +architecture arqmultisteps of multisteps is�        '      entity multisteps is5��              
          0       
              �              
          �       
              �       !       
                
              5�_�                    �   J    ����                                                                                                                                                                                                                                                                                                                            �   J       �   J          J    fYJ    �   �   �  '      ^        inst7: somador_v0 port map (a => bout, b => x"bb67ae85",  soma => haso(63 downto 32));   ^        inst8: somador_v0 port map (a => cout, b => x"3c6ef372",  soma => haso(95 downto 64));   _        inst9: somador_v0 port map (a => dout, b => x"a54ff53a",  soma => haso(127 downto 96));�   �   �  '      ]        inst6: somador_v0 port map (a => aout, b => x"6a09e667",  soma => haso(31 downto 0));5��    �   J                  �                     �    �   J                  ^                     �    �   J                  �                     �    �   J                                       5�_�                    2       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   1   2          Ksignal s1, s2, s3, s4, sa, sb, sc, sd, sW, se, sf: bit_vector(31 downto 0);5��    1                      �      L               5�_�                    4       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   3   4          signal step: integer; 5��    3                      �                     5�_�                    3   7    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   2   4  %      Wsignal aout, bout, cout, dout, eout, fout, gout, hout, kpwout: bit_vector(31 downto 0);5��    2   7                  `                     5�_�                    3   5    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   2   4  %      Qsignal aout, bout, cout, dout, eout, fout, gout, hout, : bit_vector(31 downto 0);5��    2   5                  ^                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �          &    soma : out bit_vector(31 downto 0)�   �   �          a        inst13: somador_v0 port map (a => hout, b => x"5be0cd19",  soma => haso(255 downto 224));�   �   �          a        inst12: somador_v0 port map (a => gout, b => x"1f83d9ab",  soma => haso(223 downto 192));�   �   �          a        inst11: somador_v0 port map (a => fout, b => x"9b05688c",  soma => haso(191 downto 160));�   �   �          a        inst10: somador_v0 port map (a => eout, b => x"510e527f",  soma => haso(159 downto 128));�   �   �          `        inst9: somador_v0 port map (a => dout, b => x"a54ff53a",  soma =>  haso(127 downto 96));�   �   �          _        inst8: somador_v0 port map (a => cout, b => x"3c6ef372",  soma =>  haso(95 downto 64));�   �   �          _        inst7: somador_v0 port map (a => bout, b => x"bb67ae85",  soma =>  haso(63 downto 32));�   �   �          ^        inst6: somador_v0 port map (a => aout, b => x"6a09e667",  soma =>  haso(31 downto 0));�   �   �          $                        hin <= hout;�   �   �          $                        gin <= gout;�   �   �          $                        fin <= fout;�   �   �          $                        ein <= eout;�   �   �          $                        din <= dout;�   �   �          $                        cin <= cout;�   �   �          $                        bin <= bout;�   �   �          $                        ain <= aout;�   �   �          t        inststep : stepfun port map (ain,bin,cin,din,ein,fin,gin,hin,kpwin,aout,bout,cout,dout,eout,fout,gout,hout);�   2   4          Osignal aout, bout, cout, dout, eout, fout, gout, hout: bit_vector(31 downto 0);�   (   *          &        q: out bit_vector(31 downto 0)�   !   #          &        q: out bit_vector(31 downto 0)�                &    soma : out bit_vector(31 downto 0)�                7  ao,bo,co,do,eo,fo,go,ho: out bit_vector (31 downto 0)�      
                  done : out bit�      	  %      ,        haso : out bit_vector(255 downto 0);5��                        �                     �                        �                     �                        �                    �                        7                    �    !                    �                    �    (                    A                    �    2                    7                    �    2                    >                    �    2                    E                    �    2                    L                    �    2   $                 S                    �    2   +                 Z                    �    2   2                 a                    �    2   9                 h                    �    �   L                 �                    �    �   R                 �                    �    �   X                 �                    �    �   ^                 �                    �    �   d                 �                    �    �   j                 �                    �    �   p                 �                    �    �   v                 �                    �    �                     �                    �    �                                         �    �                     <                    �    �                     b                    �    �                     �                    �    �                     �                    �    �                     �                    �    �                     �                    �    �   *                 �                    �    �   *                 �                    �    �   *                 S                    �    �   *                 �                    �    �   +                                     �    �   +                 z                    �    �   +                 �                    �    �   +                 @                    �    �                    �                    5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �  %      '    soma : _out bit_vector(31 downto 0)5��    �                     �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�      �      	  %      -        haso : _out bit_vector(255 downto 0);5��                         �                      5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                             f�     �      
  %              done : _out bit5��                         �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�     �        %      8  ao,bo,co,do,eo,fo,go,ho: _out bit_vector (31 downto 0)5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�     �        %      '    soma : _out bit_vector(31 downto 0)5��                         4                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�     �        %      &    soma : out bit_vector(31 downto 0)5��                        -                    5�_�                   %       ����                                                                                                                                                                                                                                                                                                                                                             f�     �  $              end somador_v0arch;5��    $                   Y'                    �    $                    \'                     �    $                    ['                     �    $                    Z'                     �    $                
   Y'             
       5�_�                    �       ����                                                                                                                                                                                                                                                                                                                           #          �          V       f�&     �   �   �       E   #signal c : bit_vector(31 downto 0);       begin           c(0)  <= '0';       c(1)  <= a(0) and b(0);   ;    c(2)  <= (a(1) and b(1)) or (c(1) and (a(1) xor b(1)));   ;    c(3)  <= (a(2) and b(2)) or (c(2) and (a(2) xor b(2)));   ;    c(4)  <= (a(3) and b(3)) or (c(3) and (a(3) xor b(3)));   ;    c(5)  <= (a(4) and b(4)) or (c(4) and (a(4) xor b(4)));   ;    c(6)  <= (a(5) and b(5)) or (c(5) and (a(5) xor b(5)));   ;    c(7)  <= (a(6) and b(6)) or (c(6) and (a(6) xor b(6)));   ;    c(8)  <= (a(7) and b(7)) or (c(7) and (a(7) xor b(7)));   ;    c(9)  <= (a(8) and b(8)) or (c(8) and (a(8) xor b(8)));   ;    c(10) <= (a(9) and b(9)) or (c(9) and (a(9) xor b(9)));   @    c(11) <= (a(10) and b(10)) or (c(10) and (a(10) xor b(10)));   @    c(12) <= (a(11) and b(11)) or (c(11) and (a(11) xor b(11)));   @    c(13) <= (a(12) and b(12)) or (c(12) and (a(12) xor b(12)));   @    c(14) <= (a(13) and b(13)) or (c(13) and (a(13) xor b(13)));   @    c(15) <= (a(14) and b(14)) or (c(14) and (a(14) xor b(14)));   @    c(16) <= (a(15) and b(15)) or (c(15) and (a(15) xor b(15)));   @    c(17) <= (a(16) and b(16)) or (c(16) and (a(16) xor b(16)));   @    c(18) <= (a(17) and b(17)) or (c(17) and (a(17) xor b(17)));   @    c(19) <= (a(18) and b(18)) or (c(18) and (a(18) xor b(18)));   @    c(20) <= (a(19) and b(19)) or (c(19) and (a(19) xor b(19)));   @    c(21) <= (a(20) and b(20)) or (c(20) and (a(20) xor b(20)));   @    c(22) <= (a(21) and b(21)) or (c(21) and (a(21) xor b(21)));   @    c(23) <= (a(22) and b(22)) or (c(22) and (a(22) xor b(22)));   @    c(24) <= (a(23) and b(23)) or (c(23) and (a(23) xor b(23)));   @    c(25) <= (a(24) and b(24)) or (c(24) and (a(24) xor b(24)));   @    c(26) <= (a(25) and b(25)) or (c(25) and (a(25) xor b(25)));   @    c(27) <= (a(26) and b(26)) or (c(26) and (a(26) xor b(26)));   @    c(28) <= (a(27) and b(27)) or (c(27) and (a(27) xor b(27)));   @    c(29) <= (a(28) and b(28)) or (c(28) and (a(28) xor b(28)));   @    c(30) <= (a(29) and b(29)) or (c(29) and (a(29) xor b(29)));   @    c(31) <= (a(30) and b(30)) or (c(30) and (a(30) xor b(30)));             soma(0)  <= a(0) xor b(0);   '    soma(1)  <= a(1) xor b(1) xor c(1);   '    soma(2)  <= a(2) xor b(2) xor c(2);   '    soma(3)  <= a(3) xor b(3) xor c(3);   '    soma(4)  <= a(4) xor b(4) xor c(4);   '    soma(5)  <= a(5) xor b(5) xor c(5);   '    soma(6)  <= a(6) xor b(6) xor c(6);   '    soma(7)  <= a(7) xor b(7) xor c(7);   '    soma(8)  <= a(8) xor b(8) xor c(8);   '    soma(9)  <= a(9) xor b(9) xor c(9);   *    soma(10) <= a(10) xor b(10) xor c(10);   *    soma(11) <= a(11) xor b(11) xor c(11);   *    soma(12) <= a(12) xor b(12) xor c(12);   *    soma(13) <= a(13) xor b(13) xor c(13);   *    soma(14) <= a(14) xor b(14) xor c(14);   *    soma(15) <= a(15) xor b(15) xor c(15);   *    soma(16) <= a(16) xor b(16) xor c(16);   *    soma(17) <= a(17) xor b(17) xor c(17);   *    soma(18) <= a(18) xor b(18) xor c(18);   *    soma(19) <= a(19) xor b(19) xor c(19);   *    soma(20) <= a(20) xor b(20) xor c(20);   *    soma(21) <= a(21) xor b(21) xor c(21);   *    soma(22) <= a(22) xor b(22) xor c(22);   *    soma(23) <= a(23) xor b(23) xor c(23);   *    soma(24) <= a(24) xor b(24) xor c(24);   *    soma(25) <= a(25) xor b(25) xor c(25);   *    soma(26) <= a(26) xor b(26) xor c(26);   *    soma(27) <= a(27) xor b(27) xor c(27);   *    soma(28) <= a(28) xor b(28) xor c(28);   *    soma(29) <= a(29) xor b(29) xor c(29);   *    soma(30) <= a(30) xor b(30) xor c(30);   *    soma(31) <= a(31) xor b(31) xor c(31);5��    �       E               I                    5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�(     �   �   �   �      ,architecture somador_v0arch of somador_v0 is5��    �                 
   )             
       5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�+     �   �   �   �      (architecture behavioral of somador_v0 is5��    �          
       	   7      
       	       5�_�                    �   #    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�?     �   �   �   �          �   �   �   �    �   �   �   �    5��    �                      D                     �    �                      D                     �    �                      D                     �    �                      D                    5�_�      !               �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�B    �   �   �           5��    �                      Y                     5�_�       "           !   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�w     �   �   �   �      end somador_v0;5��    �          
       	         
       	       5�_�   !   #           "   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�{     �   �   �   �      entity somador_v0 is5��    �          
       	   �      
       	       5�_�   "   $           #   �   C    ����                                                                                                                                                                                                                                                                                                                            �   C       �   C          C    f��     �   �   �   �      `        inst7: somador_v0 port map (a => b_out, b => x"bb67ae85",  soma =>  haso(63 downto 32));   `        inst8: somador_v0 port map (a => c_out, b => x"3c6ef372",  soma =>  haso(95 downto 64));   a        inst9: somador_v0 port map (a => d_out, b => x"a54ff53a",  soma =>  haso(127 downto 96));�   �   �   �      _        inst6: somador_v0 port map (a => a_out, b => x"6a09e667",  soma =>  haso(31 downto 0));5��    �   C                  �                     �    �   C                                       �    �   C                  g                     �    �   C                  �                     5�_�   #   %           $   �   E    ����                                                                                                                                                                                                                                                                                                                            �   E       �   G          G    f��     �   �   �   �      `        inst6: somador_v0 port map (a => a_out, b => x"6a09e667",   soma =>  haso(31 downto 0));   a        inst7: somador_v0 port map (a => b_out, b => x"bb67ae85",   soma =>  haso(63 downto 32));   a        inst8: somador_v0 port map (a => c_out, b => x"3c6ef372",   soma =>  haso(95 downto 64));   b        inst9: somador_v0 port map (a => d_out, b => x"a54ff53a",   soma =>  haso(127 downto 96));   b        inst10: somador_v0 port map (a => e_out, b => x"510e527f",  soma => haso(159 downto 128));   b        inst11: somador_v0 port map (a => f_out, b => x"9b05688c",  soma => haso(191 downto 160));   b        inst12: somador_v0 port map (a => g_out, b => x"1f83d9ab",  soma => haso(223 downto 192));   b        inst13: somador_v0 port map (a => h_out, b => x"5be0cd19",  soma => haso(255 downto 224));5��    �   E                  �                     �    �   E                                       �    �   E                  c                     �    �   E                  �                     �    �   E                  "                     �    �   E                  �                     �    �   E                  �                     �    �   E                  B                     5�_�   $   &           %   )       ����                                                                                                                                                                                                                                                                                                                            �   E       �   G          G    f��     �   (   *   �      '        q: _out bit_vector(31 downto 0)5��    (                     :                     5�_�   %   '           &   �   8    ����                                                                                                                                                                                                                                                                                                                            �   E       �   G          G    f��     �   �   �   �      H        	sum: somador_v0 port map(a => waux, b => kaux, soma => kpwaux);5��    �   8                 �                    5�_�   &   (           '   "       ����                                                                                                                                                                                                                                                                                                                            �   E       �   G          G    f��    �   !   #   �      '        q: _out bit_vector(31 downto 0)5��    !                     �                     5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                             f��     �         �      entity multisteps_v0 is5��                         :                      5�_�   (   *           )          ����                                                                                                                                                                                                                                                                                                                                                             f��     �         �      entity multistepsv0 is5��                         :                      5�_�   )   +           *          ����                                                                                                                                                                                                                                                                                                                                                             f��     �         �      entity multisteps0 is5��                         :                      5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                                             f��     �         �      1architecture arqmultisteps_v0 of multisteps_v0 is5��                        �                     �                     
   �              
       �              
          �       
              �                     
   �              
       5�_�   +   -           ,      %    ����                                                                                                                                                                                                                                                                                                                                                             f��     �         �      +architecture behavioral of multisteps_v0 is5��       %                                       5�_�   ,   .           -      %    ����                                                                                                                                                                                                                                                                                                                                                             f��     �         �      *architecture behavioral of multistepsv0 is5��       %                                       5�_�   -   /           .      %    ����                                                                                                                                                                                                                                                                                                                                                             f��     �         �      )architecture behavioral of multisteps0 is5��       %                                       5�_�   .   0           /   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      +        r(i) <= A(i) xor B(i) xor carry(i);5��    �                    z                    5�_�   /   1           0   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      &    soma : out bit_vector(31 downto 0)5��    �                    �                    5�_�   0               1   �       ����                                                                                                                                                                                                                                                                                                                                                             f��    �   �   �   �      +    r(31) <= A(31) xor B(31) xor carry(31);5��    �                                        5�_�                    �   #    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f�8     �   �   �   �    �   �   �   �      1architecture behavioral of somador32somador_v0 is5��    �   $               
   @              
       5�_�   	       
                 ����                                                                                                                                                                                                                                                                                                                            �   G       �   G       V   G    f6�     �        '      component somador_v0 is�   �   �          4        	inst3: somador_v0 port map(y1, W(i-7), y3);�   �   �          0        	inst4: somador_v0 port map(y3, y2, y4);�   �   �          5        	inst5: somador_v0 port map(y4, W(i-16), y5);�   �   �          H        	sum: somador_v0 port map(a => waux, b => kaux, soma => kpwaux);�   �   �          ]        inst6: somador_v0 port map (a => aout, b => x"6a09e667",  soma => haso(31 downto 0));�   �   �          ^        inst7: somador_v0 port map (a => bout, b => x"bb67ae85",  soma => haso(63 downto 32));�   �   �          ^        inst8: somador_v0 port map (a => cout, b => x"3c6ef372",  soma => haso(95 downto 64));�   �   �          _        inst9: somador_v0 port map (a => dout, b => x"a54ff53a",  soma => haso(127 downto 96));�   �   �          a        inst10: somador_v0 port map (a => eout, b => x"510e527f",  soma => haso(159 downto 128));�   �   �          a        inst11: somador_v0 port map (a => fout, b => x"9b05688c",  soma => haso(191 downto 160));�   �   �          a        inst12: somador_v0 port map (a => gout, b => x"1f83d9ab",  soma => haso(223 downto 192));�   �   �          a        inst13: somador_v0 port map (a => hout, b => x"5be0cd19",  soma => haso(255 downto 224));�   �   �          --somador_v0�   �   �          entity somador_v0 is�   �   �          end somador_v0;�   �   �          )architecture somador_v0arch of somador is�  &  (          end somador_v0arch;5��       
              
   �             
       �    �                 
   �             
       �    �                 
   �             
       �    �                 
                
       �    �                 
                
       �    �                 
   �             
       �    �                 
                
       �    �                 
   x             
       �    �                 
   �             
       �    �                 
   8             
       �    �                 
   �             
       �    �                 
   �             
       �    �                 
   ^             
       �    �                 
   �             
       �    �                 
   �             
       �    �                 
   N             
       �    �                 
   h             
       �    &                
   �'             
       5�_�   	              
   �       ����                                                                                                                                                                                                                                                                                                                            �   G       �   G       V   G    f6~     �   �   �  '      entity somadorr is5��    �                     �                     5��