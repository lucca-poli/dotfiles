Vim�UnDo� �oXp�x����S�9i�[>��m�%�uAy���   N                 	       	   	   	    f�    _�                     	       ����                                                                                                                                                                                                                                                                                                                                                             f��     �      
   V      end serial_out_tb;5��                         �                      5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                             f�      �      
   V      end ;5��                         �                      5�_�                    	        ����                                                                                                                                                                                                                                                                                                                                                             f�    �      	   V      entity serial_out_tb is   end;�      
   V      end;5��                         �                      �                         �                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f�     �                 5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�     �                 -- Testbench5��                                                  5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�     �                use IEEE.STD_LOGIC_1164.ALL;   use IEEE.STD_LOGIC_ARITH.ALL;5��                                 ;               5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�     �                 use IEEE.STD_LOGIC_UNSIGNED.ALL;5��                                 !               5�_�      	                      ����                                                                                                                                                                                                                                                                                                                                                             f�     �                 library IEEE;5��                                                  5�_�                  	           ����                                                                                                                                                                                                                                                                                                                                                             f�    �                  5��                                                  5��