Vim�UnDo� ��l�y�.�9r��b���2�Y���3�z>  �   $architecture sha256_arch of exp6 is   �                          fC�    _�                            ����                                                                                                                                                                                                                                                                                                                                       X           V        fC�l    �                  5��                                                  5�_�                   �       ����                                                                                                                                                                                                                                                                                                                                                             fC��     �  �  �  �      entity exp6 is port (5��    �                   ҁ                    5�_�                   �       ����                                                                                                                                                                                                                                                                                                                                                             fC�     �  �  �  �      	end exp6;5��    �                   6�                    5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             fC�    �  �  �  �      $architecture sha256_arch of exp6 is 5��    �                   [�                    �    �                    ]�                     �    �                    \�                     �    �                   [�                    �    �                   [�                    �    �                   [�                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                       V           V        fC�l     �              5��                                 �               5�_�                            ����                                                                                                                                                                                                                                                                                                                                       S           V        fC�m     �              5��                                 Y               5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        fC�s     �      T        5��           R                      �              5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        fC�v     �              5��                                                5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        fC�w     �               5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                                       >           V        fC�x     �               5��                                   �               5�_�      	                      ����                                                                                                                                                                                                                                                                                                                                                   V        fC��     �       ?        5��            >                                     5�_�      
           	           ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �       !        5��                                    �              5�_�   	              
           ����                                                                                                                                                                                                                                                                                                                                                V       fC��    �               5��                                                  5�_�   
                         ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �               5��                                   j              5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        fC�     �              5��                                 T              5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        fC�     �               5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        fC�     �               5��                                                  5�_�                     J       ����                                                                                                                                                                                                                                                                                                                                                  V        fC�X     �   I   K  �      U	generic(n : integer := 7); --indica o tamanho do contador(7) (bit de parada no bit7)5��    I                     �                     5�_�                             ����                                                                                                                                                                                                                                                                                                                                                  V        fC�a     �      Y        5��           T                     �              5��