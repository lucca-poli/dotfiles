Vim�UnDo� �]r�=��w�Aq�Op����k�@�JTF�����   H   entity maj_tb is end;                              e�=m    _�                             ����                                                                                                                                                                                                                                                                                                                                                             e�=]     �                   �               5��                    G                       �      5�_�                             ����                                                                                                                                                                                                                                                                                                                                                             e�=l    �                >        file tb_file : text open read_mode is "cases/maj.dat";�                    dut: maj�      
              component maj�                architecture dut of maj_tb is�         H      entity maj_tb is end;5��                        D                     �                        i                     �                        �                     �       	                 �                    �       5                 �                    5��