Vim�UnDo� �9&	Z��(9��?���sZdV�s)/	v��979   �   !    component interface_hcsr04 is   0                           fs�    _�                      0        ����                                                                                                                                                                                                                                                                                                                                                             fs�    �   n   p              sensor: interface_hcsr04�   <   >           	end component interface_hcsr04;�   /   1   �      !    component interface_hcsr04 is5��    /                    �                    �    <                    -                    �    n                    |                    5��