Vim�UnDo� ����Y�ie
�85�C�8��LT}%��   D   =            " B=" & integer'image(to_integer(signed(y))) &LF&   7   4      1       1   1   1    e�"    _�                             ����                                                                                                                                                                                                                                                                                                                                                             e�!A     �   A   C          <        assert false report "EOT ch function" severity note;�   "   $          <        assert false report "BOT ch function" severity note;�                "        variable space: character;�                =        file tb_file : text open read_mode is "cases/ch.dat";�                    dut: ch�                     -- Signals for the testbench�      
              component ch�                architecture dut of ch_tb is�         G      entity ch_tb is end;5��                        D                     �                        Z                     �                        �                     �                        u                    �       	                                     �       5                 �                    �                        �                    �    "   !                 ~                    �    A   !                 D                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 v       e�!b     �         G      !arsomadoritecture dut of ch_tb is�         G    5��                         X                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 v       e�!f     �         G      architecture dut of ch_tb is5��                        l                     �                         n                      �                         m                      �                        l                     �                     
   l              
       �              
       
   l       
       
       �              
          l       
              �                     
   l              
       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 v       e�!l     �         G      '        variable space: somadoraracter;5��                        �                    �                         �                     �                        �                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            .          /          V       e�!�     �          G      :        variable Xv, Yv, Zv, res: bit_vector(31 downto 0);5��                                              5�_�                           ����                                                                                                                                                                                                                                                                                                                            .          /          V       e�!�     �          G      8        variable Xv, Yv, , res: bit_vector(31 downto 0);5��                                              5�_�                           ����                                                                                                                                                                                                                                                                                                                            .          /          V       e�!�     �          G      6        variable Xv, Yv, res: bit_vector(31 downto 0);5��                                            5�_�                           ����                                                                                                                                                                                                                                                                                                                            .          /          V       e�!�     �          G      6        variable Av, Yv, res: bit_vector(31 downto 0);5��                                            5�_�                    )       ����                                                                                                                                                                                                                                                                                                                            .          /          V       e�!�     �   (   *   G                  read(tb_line, Xv);5��    (                                        5�_�                    )       ����                                                                                                                                                                                                                                                                                                                            .          /          V       e�!�     �   (   *   G                  read(tb_line, av);5��    (                                        5�_�                    ,       ����                                                                                                                                                                                                                                                                                                                            .          /          V       e�!�     �   +   -   G                  read(tb_line, Yv);5��    +                    s                    5�_�                    .       ����                                                                                                                                                                                                                                                                                                                            .          /          V       e�!�     �   -   .          !            read(tb_line, space);               read(tb_line, Zv);5��    -                      �      A               5�_�                    .       ����                                                                                                                                                                                                                                                                                                                            .          .          V       e�!�     �   -   .                      z <= Zv;5��    -                      �                     5�_�                    *       ����                                                                                                                                                                                                                                                                                                                            .          .          V       e�!�     �   )   +   D                  x <= Xv;5��    )                    3                    5�_�                    -       ����                                                                                                                                                                                                                                                                                                                            .          .          V       e�!�     �   ,   .   D                  y <= Yv;5��    ,                    �                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       e�!�     �   
      B    �         B    �   
             0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)5��    
                      �       \               �    
                      �               x       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �         E      '        B : in bit_vector(31 downto 0);   '        S : out bit_vector(31 downto 0)�   
      E      '        A : in bit_vector(31 downto 0);5��    
                     �                      �                                              �                         <                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �         E      6        port map (x => x, y => y, z => z, q => saida);5��                        E                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �         E      6        port map (A => x, y => y, z => z, q => saida);5��                        J                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �         E      6        port map (A => A, y => y, z => z, q => saida);5��                        M                    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �         E      6        port map (A => A, A => y, z => z, q => saida);5��                        R                    5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �         E      6        port map (A => A, A => A, z => z, q => saida);5��                        R                    5�_�       "           !          ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �         E      6        port map (A => A, A => B, z => z, q => saida);5��                        M                    5�_�   !   #           "           ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �         E      6        port map (A => A, B => B, z => z, q => saida);5��                          S                     5�_�   "   $           #      "    ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �         E      .        port map (A => A, B => B, q => saida);5��       "                 U                    5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �         E      -    signal x, y, z : bit_vector(31 downto 0);5��                         �                     5�_�   $   &           %          ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �         E      +    signal x, y, : bit_vector(31 downto 0);5��                         �                     5�_�   %   '           &          ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �         E      *    signal x, y : bit_vector(31 downto 0);5��                        �                    5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �         E      *    signal x, B : bit_vector(31 downto 0);5��                        �                    5�_�   '   )           (   +       ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �   *   ,   E                  x <= Av;5��    *                    K                    5�_�   (   *           )   .       ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �   -   /   E                  y <= Bv;5��    -                    �                    5�_�   )   +           *   8       ����                                                                                                                                                                                                                                                                                                                                                       e�!�     �   7   8          =            " Z=" & integer'image(to_integer(signed(z))) &LF&5��    7                      �      >               5�_�   *   ,           +   8       ����                                                                                                                                                                                                                                                                                                                                                       e�"     �   7   9   D      J            " Computed Q=" & integer'image(to_integer(signed(saida))) &LF&5��    7                    �                    5�_�   +   -           ,   9       ����                                                                                                                                                                                                                                                                                                                                                       e�"     �   8   :   D      C            " Expected Q=" & integer'image(to_integer(signed(res)))5��    8                    .                    5�_�   ,   .           -   6       ����                                                                                                                                                                                                                                                                                                                                                       e�"	     �   5   7   D      =            " X=" & integer'image(to_integer(signed(x))) &LF&5��    5                    ^                    5�_�   -   /           .   7       ����                                                                                                                                                                                                                                                                                                                                                       e�"     �   6   8   D      =            " Y=" & integer'image(to_integer(signed(y))) &LF&5��    6                    �                    5�_�   .   0           /   6   4    ����                                                                                                                                                                                                                                                                                                                                                       e�"     �   5   7   D      =            " A=" & integer'image(to_integer(signed(x))) &LF&5��    5   4                 �                    5�_�   /   1           0   7   4    ����                                                                                                                                                                                                                                                                                                                                                       e�"     �   6   8   D      =            " B=" & integer'image(to_integer(signed(y))) &LF&5��    6   4                 �                    5�_�   0               1   7   4    ����                                                                                                                                                                                                                                                                                                                                                       e�"    �   6   8   D      =            " B=" & integer'image(to_integer(signed(A))) &LF&5��    6   4                 �                    5�_�                         ����                                                                                                                                                                                                                                                                                                                                                             e�!M     �         G       aromadoritecture dut of ch_tb is5��                         Z                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�!N     �         G      armadoritecture dut of ch_tb is5��                         Z                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�!N     �         G      aradoritecture dut of ch_tb is5��                         Z                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�!N     �         G      ardoritecture dut of ch_tb is5��                         Z                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�!N     �         G      aroritecture dut of ch_tb is5��                         Z                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�!N     �         G      arritecture dut of ch_tb is5��                         Z                      5�_�          	                 ����                                                                                                                                                                                                                                                                                                                                                             e�!S     �         G      arcitecture dut of ch_tb is5��                        Z                     5�_�      
          	          ����                                                                                                                                                                                                                                                                                                                                                             e�!N     �         G      aritecture dut of ch_tb is5��                         Z                      5�_�   	               
          ����                                                                                                                                                                                                                                                                                                                                                             e�!O     �         G      artecture dut of ch_tb is5��                         Z                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             e�!H     �         G      arch dut of ch_tb is5��                         X                     5��