Vim�UnDo� W.����k����@ȩ�yG�):�o)�v��g   �                  I       I   I   I    fB��   
 _�                     W        ����                                                                                                                                                                                                                                                                                                                            ;          W          V       f:s�     �   W               �   W            5��    W                      �                     �    W                      �                     5�_�                    X       ����                                                                                                                                                                                                                                                                                                                            ;          W          V       f:s�     �   W              p5��    W                      �                     5�_�                    X        ����                                                                                                                                                                                                                                                                                                                            ;          W          V       f:s�     �   X            �   X            5��    X                      �              x      5�_�                    \       ����                                                                                                                                                                                                                                                                                                                            ;          W          V       f:s�     �   [   ]   u      entity shift_reg512 is5��    [                    5                    5�_�                    o       ����                                                                                                                                                                                                                                                                                                                            ;          W          V       f:t�     �   n   p   u      2            vector <= vector(479 downto 0) & data;5��    n                    	                    5�_�                    _       ����                                                                                                                                                                                                                                                                                                                            ;          W          V       f:t�     �   ^   `   u      )        data: in bit_vector(31 downto 0);5��    ^                    �                    5�_�                    c       ����                                                                                                                                                                                                                                                                                                                            ;          W          V       f:t�     �   b   d   u      end entity shift_reg512;5��    b   
                  �                     5�_�      	              e   #    ����                                                                                                                                                                                                                                                                                                                            ;          W          V       f:t�    �   d   f   u      (architecture Behavior of shift_reg512 is5��    d   #                                       �    d   "                                     �    d   #                                       �    d   "                                       �    d   !                                       �    d                                           �    d                                          �    d                                          �    d                                          �    d                                          �    d                                          �    d                                          �    d                                        �    d                 	                	       �    d          	                	              5�_�      
           	   `       ����                                                                                                                                                                                                                                                                                                                            ;          W          V       f:�#     �   _   `          '        d: in bit_vector(511 downto 0);5��    _                      �      (               5�_�   	              
   l       ����                                                                                                                                                                                                                                                                                                                            ;          W          V       f:�'     �   k   m   t                  vector <= d;5��    k                     �                     5�_�   
                 l       ����                                                                                                                                                                                                                                                                                                                            ;          W          V       f:�(     �   k   m   t                  vector <= ;5��    k                     �                     5�_�                    l       ����                                                                                                                                                                                                                                                                                                                            ;          W          V       f:�)    �   k   m   t                  vector <= ();5��    k                     �                     �    k                    �                    �    k                    �                    �    k                    �                    �    k                    �                    5�_�                            ����                                                                                                                                                                                                                                                                                                                                      9          V       f:�5     �         t    5��                          =                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                      :          V       f:�6     �      :   u    �         u    5��                          >              D      5�_�                    !   
    ����                                                                                                                                                                                                                                                                                                                            ;          V          V       f:�<     �       "   �      entity reg32 is5��        
                 q                    5�_�                    (       ����                                                                                                                                                                                                                                                                                                                            ;          V          V       f:�J     �   '   )   �      end entity reg32;5��    '                     /                     5�_�                    (       ����                                                                                                                                                                                                                                                                                                                            ;          V          V       f:�K     �   '   )   �      end entity ;5��    '   
                  .                     5�_�                    $       ����                                                                                                                                                                                                                                                                                                                            ;          V          V       f:�v     �   #   $          )        init: in bit_vector(31 downto 0);5��    #                      �      *               5�_�                    0       ����                                                                                                                                                                                                                                                                                                                            :          U          V       f:�y     �   /   1   �                  value <= init;5��    /                     �                     5�_�                    0       ����                                                                                                                                                                                                                                                                                                                            :          U          V       f:�z     �   /   1   �                  value <= ;5��    /                     �                     5�_�                    0       ����                                                                                                                                                                                                                                                                                                                            :          U          V       f:�{     �   /   1   �                  value <= "";5��    /                     �                     5�_�                    0       ����                                                                                                                                                                                                                                                                                                                            :          U          V       f:�{     �   /   1   �                  value <= ;5��    /                     �                     5�_�                    0       ����                                                                                                                                                                                                                                                                                                                            :          U          V       f:�|     �   /   1   �                  value <= ();5��    /                     �                     �    /                    �                    �    /                    �                    �    /                    �                    �    /                    �                    5�_�                    )       ����                                                                                                                                                                                                                                                                                                                            :          U          V       f:��     �   (   *   �      !architecture Behavior of reg32 is5��    (                    #                    5�_�                    *       ����                                                                                                                                                                                                                                                                                                                            :          U          V       f:��     �   )   +   �      *    signal value: bit_vector(31 downto 0);5��    )                    G                    5�_�                    $       ����                                                                                                                                                                                                                                                                                                                            :          U          V       f:��     �   #   %   �      &        d: in bit_vector(31 downto 0);5��    #                    �                    5�_�                    %       ����                                                                                                                                                                                                                                                                                                                            :          U          V       f:��    �   $   &   �      &        q: out bit_vector(31 downto 0)5��    $                    �                    5�_�                            ����                                                                                                                                                                                                                                                                                                                                      9           V       f:��    �                library IEEE;   use IEEE.NUMERIC_BIT.all;       entity reg512 is   
    port (   !        rst, clk, enable: in bit;   '        d: in bit_vector(511 downto 0);   '        q: out bit_vector(511 downto 0)       );   end entity;       "architecture Behavior of reg512 is   +    signal value: bit_vector(511 downto 0);   begin              process(rst, clk)   	    begin           if rst = '1' then   %            value <= (others => '0');   4        elsif rising_edge(clk) and enable = '1' then               value <= D;           end if;       end process;           q <= value;          end architecture Behavior;    5��                          >      %              5�_�                    W        ����                                                                                                                                                                                                                                                                                                                            Y           t           V        f;g�     �   W   Y   t    5��    W                      �                     5�_�                    X        ����                                                                                                                                                                                                                                                                                                                            Z           u           V        f;g�     �   X   u   u    �   X   Y   u    5��    X                      �              T      5�_�                     \       ����                                                                                                                                                                                                                                                                                                                            v           �           V        f;g�     �   [   ]   �      entity shift_reg_byte is5��    [                     :                     5�_�      !               _       ����                                                                                                                                                                                                                                                                                                                            v           �           V        f;g�     �   ^   `   �      (        data: in bit_vector(7 downto 0);5��    ^                    �                    5�_�       "           !   _       ����                                                                                                                                                                                                                                                                                                                            v           �           V        f;g�     �   ^   `   �      *        data: in bit_vector(255 downto 0);5��    ^                    w                    5�_�   !   #           "   `       ����                                                                                                                                                                                                                                                                                                                            v           �           V        f;g�     �   _   a   �      '        q: out bit_vector(511 downto 0)5��    _                    �                    5�_�   "   $           #   d   '    ����                                                                                                                                                                                                                                                                                                                            v           �           V        f;g�     �   c   e   �      *architecture Behavior of shift_reg_byte is5��    c   '                  �                     5�_�   #   %           $   e       ����                                                                                                                                                                                                                                                                                                                            v           �           V        f;h     �   d   f   �      ,   signal vector: bit_vector(511 downto 0); 5��    d                                        5�_�   $   &           %   n       ����                                                                                                                                                                                                                                                                                                                            v           �           V        f;h     �   m   o   �      2            vector <= vector(503 downto 0) & data;5��    m                    �                    5�_�   %   '           &   m       ����                                                                                                                                                                                                                                                                                                                            v           �           V        f;h�     �   l   n   �      4        elsif rising_edge(clk) and enable = '1' then5��    l                     �                     5�_�   &   (           '   m       ����                                                                                                                                                                                                                                                                                                                            v           �           V        f;h�     �   l   n   �      0        elsif rising_edge(clk) enable = '1' then5��    l                     �                     5�_�   '   )           (   m       ����                                                                                                                                                                                                                                                                                                                            v           �           V        f;h�     �   l   n   �      )        elsif rising_edge(clk) = '1' then5��    l                     �                     5�_�   (   *           )   m       ����                                                                                                                                                                                                                                                                                                                            v           �           V        f;h�     �   l   n   �      '        elsif rising_edge(clk) '1' then5��    l                     �                     5�_�   )   +           *   m       ����                                                                                                                                                                                                                                                                                                                            v           �           V        f;h�     �   l   n   �      &        elsif rising_edge(clk) 1' then5��    l                     �                     5�_�   *   ,           +   m       ����                                                                                                                                                                                                                                                                                                                            v           �           V        f;h�     �   l   n   �      %        elsif rising_edge(clk) ' then5��    l                     �                     5�_�   +   -           ,   n       ����                                                                                                                                                                                                                                                                                                                            v           �           V        f;h�     �   m   o   �                  �   m   o   �    5��    m                      �                     �    m                     �                     �    m                     �                     �    m                     �                     �    m                    �                    �    m                    �                    �    m                 	   �             	       5�_�   ,   .           -   n       ����                                                                                                                                                                                                                                                                                                                            w           �           V        f;h�     �   m   o   �                  if enable = 5��    m                     �                     5�_�   -   /           .   n       ����                                                                                                                                                                                                                                                                                                                            w           �           V        f;h�     �   m   o   �                  if enable = ''5��    m                     �                     5�_�   .   0           /   n       ����                                                                                                                                                                                                                                                                                                                            w           �           V        f;h�     �   m   p   �                  if enable = '1'5��    m                     �                     �    m                    �                    �    m                    �                    �    m                    �                    �    m                     �                     �    n                     �                    �    n                      �                     5�_�   /   1           0   p       ����                                                                                                                                                                                                                                                                                                                            x           �           V        f;h�     �   o   p                      vector <= d;5��    o                      �                     5�_�   0   2           1   o        ����                                                                                                                                                                                                                                                                                                                            w           �           V        f;h�     �   n   p   �    �   o   p   �    5��    n                      �                     5�_�   1   3           2   o       ����                                                                                                                                                                                                                                                                                                                            x           �           V        f;h�     �   n   p   �                  vector <= d;5��    n                     �                     5�_�   2   4           3   p        ����                                                                                                                                                                                                                                                                                                                            x           �           V        f;h�     �   p   r   �                      vector�   o   r   �       5��    o                      �                     �    o                    	                    �    o                     	                     �    o                    	                     �    p                     	                    �    p                     	                     �    p                    	                    �    p                     	                     �    p                     	                     �    p                    	                    �    p                    	                    �    p                    	                    �    p                     )	                     �    p                     (	                     �    p                    '	                    �    p                    '	                    �    p                    '	                    5�_�   3   5           4   u       ����                                                                                                                                                                                                                                                                                                                            y           �           V        f;i�     �   t   v   �          q <= vector;5��    t                     _	                     5�_�   4   6           5   u       ����                                                                                                                                                                                                                                                                                                                            y           �           V        f;i�     �   t   v   �          q <= vector();5��    t                  	   `	              	       �    t                    h	                    5�_�   5   7           6   q        ����                                                                                                                                                                                                                                                                                                                            y           �           V        f;i�     �   p   r   �                       vector <= vector5��    p                      -	                     5�_�   6   8           7   q   !    ����                                                                                                                                                                                                                                                                                                                            y           �           V        f;i�     �   p   r   �      "                vector <= vector()5��    p   !                  .	                     �    p   %                 2	                    �    p   %                 2	                    �    p   %                 2	                    5�_�   7   9           8   q   .    ����                                                                                                                                                                                                                                                                                                                            y           �           V        f;i�     �   p   r   �      .                vector <= vector(247 downto 0)5��    p   .                  ;	                     5�_�   8   :           9   q   1    ����                                                                                                                                                                                                                                                                                                                            y           �           V        f;i�     �   p   r   �      1                vector <= vector(247 downto 0) & 5��    p   1                  >	                     5�_�   9   ;           :   q   2    ����                                                                                                                                                                                                                                                                                                                            y           �           V        f;i�     �   p   r   �      3                vector <= vector(247 downto 0) & ()5��    p   2                  ?	                     �    p   2                 ?	                    �    p   2                 ?	                    �    p   2                 ?	                    �    p   2                 ?	                    5�_�   :   <           ;   q   @    ����                                                                                                                                                                                                                                                                                                                            y           �           V        f;i�     �   p   r   �      @                vector <= vector(247 downto 0) & (others => '0')5��    p   @                  M	                     5�_�   ;   =           <   q   @    ����                                                                                                                                                                                                                                                                                                                            y           �           V        f;i�    �   q   s   �                      �   q   s   �    5��    q                      O	                     �    q                     _	                     �    q                     O	                    �    q                     _	                     5�_�   <   >           =   q   1    ����                                                                                                                                                                                                                                                                                                                            z           �           V        f;j�     �   p   r   �      A                vector <= vector(247 downto 0) & (others => '0');5��    p   1                  >	                     5�_�   =   ?           >   q   1    ����                                                                                                                                                                                                                                                                                                                            z           �           V        f;j�     �   p   r   �      2                vector <= vector(247 downto 0) & ;5��    p   1                  >	                     5�_�   >   @           ?   q   2    ����                                                                                                                                                                                                                                                                                                                            z           �           V        f;j�    �   p   r   �      4                vector <= vector(247 downto 0) & "";5��    p   2                  ?	                     5�_�   ?   A           @   i       ����                                                                                                                                                                                                                                                                                                                            ]   	       a          V        f;n�    �   h   j   �          process(rst, clk)5��    h                     M                     �    h                     P                     �    h                    O                    �    h                     Q                     �    h                     P                     �    h                    O                    �    h                    O                    �    h                    O                    5�_�   @   B           A   l       ����                                                                                                                                                                                                                                                                                                                            ]   	       a          V        f;s�     �   k   m   �      &            vector <= (others => '0');5��    k                    �                    5�_�   A   C           B   p       ����                                                                                                                                                                                                                                                                                                                            ]   	       a          V        f;s�     �   o   p                      else5��    o                      �                     5�_�   B   D           C   o       ����                                                                                                                                                                                                                                                                                                                            ]   	       a          V        f;s�    �   n   o                          vector <= d;5��    n                      �                     5�_�   C   E           D   !        ����                                                                                                                                                                                                                                                                                                                            !           9           V        fB��     �       =   z    �   !   "   z    �       !          entity reg32 is   
    port (   !        rst, clk, enable: in bit;   )        init: in bit_vector(31 downto 0);   &        d: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)       );   end entity reg32;       !architecture Behavior of reg32 is   *    signal value: bit_vector(31 downto 0);   begin              process(rst, clk)   	    begin           if rst = '1' then               value <= init;   4        elsif rising_edge(clk) and enable = '1' then               value <= D;           end if;       end process;           q <= value;          end architecture Behavior;5��                           g                    �                           g              D      5�_�   D   F           E           ����                                                                                                                                                                                                                                                                                                                            !           <          V        fB��     �                library IEEE;   use IEEE.NUMERIC_BIT.all;    5��                          >      )               5�_�   E   G           F   ;        ����                                                                                                                                                                                                                                                                                                                            ;          W          V       fB��     �   :   ;          library IEEE;   use IEEE.NUMERIC_BIT.all;       entity shift_reg512 is   
    port (   !        rst, clk, enable: in bit;   )        data: in bit_vector(31 downto 0);   '        d: in bit_vector(511 downto 0);   '        q: out bit_vector(511 downto 0)       );   end entity shift_reg512;       (architecture Behavior of shift_reg512 is   ,   signal vector: bit_vector(511 downto 0);        begin              process(rst, clk)   	    begin           if rst = '1' then               vector <= d;   4        elsif rising_edge(clk) and enable = '1' then   2            vector <= vector(479 downto 0) & data;           end if;       end process;           q <= vector;          end architecture Behavior;5��    :                      �      x              5�_�   F   H           G   ;        ����                                                                                                                                                                                                                                                                                                                            ;          ;          V       fB��   	 �   :   X   v    �   ;   <   v    5��    :                      �              x      5�_�   G   I           H   <        ����                                                                                                                                                                                                                                                                                                                            W           ;           V        fB��     �   :   Y   w      library IEEE;�   ;   <   w    �   ;   <          use IEEE.NUMERIC_BIT.all;       entity shift_reg512 is   
    port (   !        rst, clk, enable: in bit;   )        data: in bit_vector(31 downto 0);   '        d: in bit_vector(511 downto 0);   '        q: out bit_vector(511 downto 0)       );   end entity shift_reg512;       (architecture Behavior of shift_reg512 is   ,   signal vector: bit_vector(511 downto 0);        begin              process(rst, clk)   	    begin           if rst = '1' then               vector <= d;   4        elsif rising_edge(clk) and enable = '1' then   2            vector <= vector(479 downto 0) & data;           end if;       end process;           q <= vector;          end architecture Behavior;5��    ;                      �      j              �    :                      �                     �    :                      �              y      5�_�   H               I   X        ����                                                                                                                                                                                                                                                                                                                            Y           ;           V        fB��   
 �   W   X           5��    W                      �                     5��