Vim�UnDo� �m���z	+�YZO�.o�D������?�ԗ����   �                                   fC��    _�                            ����                                                                                                                                                                                                                                                                                                                            &                    V       f:u�     �          �    5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                            '                    V       f:u�     �       '   �    �         �    5��                    &                       �      5�_�                           ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:u�     �         �      entity counter_generic is5��                         ?                      5�_�                    	       ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:u�     �      
   �      J        clk, rst, start: in bit;                            -- Clock input5��                        �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:u�     �         �      end counter_generic;5��                        5                    5�_�                       *    ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:u�     �         �      -architecture Behavioral of counter_generic is5��       *                  h                     �       *                  h                     �       )                  g                     �       (                  f                     �       '                  e                     �       &                  d                     �       %                  c                     �       $                  b                     �       #                  a                     �       "                  `                     �       !                  _                     �                          ^                     �                         ]                     �                         \                     �                         [                     �                         Z                     �                        Y                    �                        Y                    �                        Y                    5�_�                            ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:u�     �         �      &    counting: process(clk, rst, start)5��                         �                    �       "                  �                     �       !                  �                     �                         �                    �                         �                    �                         �                    5�_�      	                     ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:v-     �         �      \            if (counter > 0 and counter < MAX_COUNT-1) or (start = '1' and counter = 0) then5��              '           �      '               5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:v.     �         �      5            if  or (start = '1' and counter = 0) then5��                         �                     5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:v/     �         �      2            if  (start = '1' and counter = 0) then5��                         �                     5�_�   
                        ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:v1     �         �      0            if(start = '1' and counter = 0) then5��                         �                     5�_�                          ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:vy     �         �      1            if (start = '1' and counter = 0) then5��                        �                    �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    �                        �                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:v~     �         �                  if enable =  then5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:v�     �         �                  if enable = '' then5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:v�     �                            end if;5��                          �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            L          '          V       f:v�     �         �                   if enable = '1' then5��                         �                     �                         �                    �                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            L          '          V       f:v�     �         �      '                elsif enable = '1' then5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            L          '          V       f:v�     �          �                      �          �    5��                          �                     �                                              �                                              �                                              �                                            �                                            �                     
                
       �                                              �                                              5�_�                           ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:v�     �          �                      done <= 5��                                              5�_�                           ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:v�     �          �                      done <= ''5��                                              5�_�                           ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:v�    �          �                      done <= '0'5��                                              5�_�                    O        ����                                                                                                                                                                                                                                                                                                                            O          o          V       fB��     �   N   n   �    �   O   P   �    �   N   O       !   library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity counter_6bit is   
    port (   C        clk, rst: in bit;                            -- Clock input           done: out bit;   O        count : out unsigned(5 downto 0)       -- 6-bit count output (64 steps)       );   end counter_6bit;       #architecture rtl of counter_6bit is   )    signal counter: unsigned(5 downto 0);       begin              counting: process(clk, rst)   	    begin           if rst = '1' then   '            counter <= (others => '0');               done <= '0';   #        elsif rising_edge(clk) then   ,            if to_integer(counter) = 63 then                   done <= '1';               else   '                counter <= counter + 1;               end if;           end if;       end process counting;           count <= counter;          end architecture rtl;5��    N       !               '                    �    N                      '              �      5�_�                    o        ����                                                                                                                                                                                                                                                                                                                            o          �          V       fB��    �   n   �   �    �   o   p   �    �   n   o          entity adder32 is   port(   &    a, b : in bit_vector(31 downto 0);   #    s : out bit_vector(31 downto 0)       );   end adder32;       %architecture behavioral of adder32 is   +    signal carry : bit_vector(31 downto 0);   begin   "    sum: for i in 0 to 30 generate   +        s(i) <= A(i) xor B(i) xor carry(i);   T        carry(i+1) <= (A(i) and B(i)) or (A(i) and carry(i)) or (B(i) and carry(i));       end generate;       +    s(31) <= A(31) xor B(31) xor carry(31);         end behavioral;5��    n                       
      �              �    n                       
              �      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        fC�Q     �          �    5��                                                  5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        fC�S     �          �    �         �    5��                                           )       5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        fC�T     �      	   �      end entity �         �      
entity  is�      	   �              �         �       �         �    5��                          )                      �                          )                      �                         +                      �                         *                      �                         )                     �                         )                     �                         )                     �                         )                     �                        0                      �                          G                       �                        G                      �                         Z                      �                      
   0               
       �                      
   d               
       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       fC�W     �         �    �      	   �      end entity components;�         �    �         �    �         �    �         �    �         �    �         �    �         �      entity components is5��              
          0       
              �              
          [       
              �                         1                      �                        \                     �       	                  2                      �                        ]                     �       
                  3                      �                        ^                     �                         4                      �                        _                     �                         5                      �                        `                     �                         6                      �                        a                     �                         N                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V        fC��    �                 library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity sampler is   
    port (   !        rst, clk, enable: in bit;       );   end entity sampler;5��                                   �               5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        fC�Q     �         �    �         �      library IEEE;   use IEEE.NUMERIC_BIT.ALL;    5��                                         )       5�_�                           ����                                                                                                                                                                                                                                                                                                                            M          (          V       f:vt     �         �      0            if start = '1' and counter = 0) then5��                         �                     5��