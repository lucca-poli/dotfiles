Vim�UnDo� \w!j�8�'�;?��R�bҘݻ͓���a:   <           %      %       %   %   %    f�f   
 _�                     ]        ����                                                                                                                                                                                                                                                                                                                            ]          o          V       f=�    �   \   ]          entity somador is   
    port (   '        A : in bit_vector(31 downto 0);   '        B : in bit_vector(31 downto 0);   '        S : out bit_vector(31 downto 0)       );   end entity somador;       %architecture behavioral of somador is   +    signal carry : bit_vector(31 downto 0);   begin   "    sum: for i in 0 to 30 generate   +        S(i) <= A(i) xor B(i) xor carry(i);   T        carry(i+1) <= (A(i) and B(i)) or (A(i) and carry(i)) or (B(i) and carry(i));       end generate;       +    S(31) <= A(31) xor B(31) xor carry(31);          end architecture behavioral;5��    \                      V
                    5�_�                            ����                                                                                                                                                                                                                                                                                                                            [           F           V        f=�    �                use IEEE.STD_LOGIC_1164.ALL;5��                                                5�_�                            ����                                                                                                                                                                                                                                                                                                                            Z           E           V        f=�     �                use IEEE.NUMERIC_STD.ALL;5��                                                5�_�                            ����                                                                                                                                                                                                                                                                                                                            Y           D           V        f=�     �                 library IEEE;5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                            X           C           V        f=�    �                  5��                                                  5�_�                   '        ����                                                                                                                                                                                                                                                                                                                                                             fm�     �   L   N          M    getA: somador port map (A => sum0Out, B => sum0Complement, S => preAOut);�   K   M          _    getSum0Complement: somador port map (A => majOut, B => majComplement, S => sum0Complement);�   J   L          G    getE: somador port map (A => di, B => majComplement, S => preEOut);�   I   K          _    getMajComplement: somador port map (A => sum1Out, B => sum1Complement, S => majComplement);�   H   J          ]    getSum1Complement: somador port map (A => chOut, B => chComplement, S => sum1Complement);�   G   I          M    getChComplement: somador port map (A => hi, B => kpw, S => chComplement);�   &   (   X          component somador is5��    &                    �                    �    G                    �                    �    H                    �                    �    I                    D                    �    J   
                 �                    �    K                    �                    �    L   
                 @	                    5�_�      	              H   :    ����                                                                                                                                                                                                                                                                                                                                                             fm�     �   G   I   X      M    getChComplement: adder32 port map (A => hi, B => kpw, S => chComplement);5��    G   :                 �                    5�_�      
           	   I   H    ����                                                                                                                                                                                                                                                                                                                                                             fm�     �   H   J   X      ]    getSum1Complement: adder32 port map (A => chOut, B => chComplement, S => sum1Complement);5��    H   H                                     5�_�   	              
   J   K    ����                                                                                                                                                                                                                                                                                                                                                             fm�     �   I   K   X      _    getMajComplement: adder32 port map (A => sum1Out, B => sum1Complement, S => majComplement);5��    I   K                 y                    5�_�   
                 K   9    ����                                                                                                                                                                                                                                                                                                                                                             fm�     �   J   L   X      G    getE: adder32 port map (A => di, B => majComplement, S => preEOut);5��    J   9                 �                    5�_�                    L   J    ����                                                                                                                                                                                                                                                                                                                                                             fm�     �   K   M   X      _    getSum0Complement: adder32 port map (A => majOut, B => majComplement, S => sum0Complement);5��    K   J                  	                    5�_�                    M   ?    ����                                                                                                                                                                                                                                                                                                                                                             fm�     �   L   N   X      M    getA: adder32 port map (A => sum0Out, B => sum0Complement, S => preAOut);5��    L   ?                 u	                    5�_�                    +       ����                                                                                                                                                                                                                                                                                                                                                             fm�    �   *   ,   X      +            S : out bit_vector(31 downto 0)5��    *                    +                    5�_�                    '        ����                                                                                                                                                                                                                                                                                                                                                             f��    �   L   N          M    getA: adder32 port map (A => sum0Out, B => sum0Complement, R => preAOut);�   K   M          _    getSum0Complement: adder32 port map (A => majOut, B => majComplement, R => sum0Complement);�   J   L          G    getE: adder32 port map (A => di, B => majComplement, R => preEOut);�   I   K          _    getMajComplement: adder32 port map (A => sum1Out, B => sum1Complement, R => majComplement);�   H   J          ]    getSum1Complement: adder32 port map (A => chOut, B => chComplement, R => sum1Complement);�   G   I          M    getChComplement: adder32 port map (A => hi, B => kpw, R => chComplement);�   &   (   X          component adder32 is5��    &                 	   �             	       �    G                 	   �             	       �    H                 	   �             	       �    I                 	   J             	       �    J   
              	   �             	       �    K                 	   �             	       �    L   
              	   L	             	       5�_�                            ����                                                                                                                                                                                                                                                                                                                                       X           V        f�[     �              X   entity stepfun is   
    port (   @    	ai, bi, ci, di, ei, fi, gi, hi: in bit_vector(31 downto 0);   (        kpw: in bit_vector(31 downto 0);   C        ao, bo, co, do, eo, fo, go, ho: out bit_vector(31 downto 0)   
        );   end stepfun;       %architecture behavioral of stepfun is   #    -- Declaração dos componentes       component ch is           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component maj is           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component sum0 is           port (   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component sum1 is           port (   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component somador32 is           port (   +            A : in bit_vector(31 downto 0);   +            B : in bit_vector(31 downto 0);   +            R : out bit_vector(31 downto 0)   
        );       end component;           -- Sinais           -- Sums complements   1    signal chComplement: bit_vector(31 downto 0);   2    signal majComplement: bit_vector(31 downto 0);   3    signal sum0Complement: bit_vector(31 downto 0);   3    signal sum1Complement: bit_vector(31 downto 0);       "    -- Crytografy funcions outputs   +    signal chOut: bit_vector(31 downto 0);    ,    signal majOut: bit_vector(31 downto 0);    -    signal sum0Out: bit_vector(31 downto 0);    -    signal sum1Out: bit_vector(31 downto 0);            -- Intermediate outputs   ,    signal preAOut: bit_vector(31 downto 0);   ,    signal preEOut: bit_vector(31 downto 0);       begin       -- Saida dos Componentes   +    getCh: ch port map (ei, fi, gi, chOut);   .    getMaj: maj port map (ai, bi, ci, majOut);   )    getSum0: sum0 port map (ai, sum0Out);   )    getSum1: sum1 port map (ei, sum1Out);       O    getChComplement: somador32 port map (A => hi, B => kpw, R => chComplement);   _    getSum1Complement: somador32 port map (A => chOut, B => chComplement, R => sum1Complement);   a    getMajComplement: somador32 port map (A => sum1Out, B => sum1Complement, R => majComplement);   I    getE: somador32 port map (A => di, B => majComplement, R => preEOut);   a    getSum0Complement: somador32 port map (A => majOut, B => majComplement, R => sum0Complement);   O    getA: somador32 port map (A => sum0Out, B => sum0Complement, R => preAOut);           ao <= preAOut;       bo <= ai;       co <= bi;       do <= ci;       eo <= preEOut;       fo <= ei;       go <= fi;       ho <= gi;   end behavioral;    5��            X                      
             5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        f�e     �                   �               5��                    X                       
      5�_�                    Y        ����                                                                                                                                                                                                                                                                                                                                                  V        f�f    �   X   Y           5��    X                      
                     5�_�                    '        ����                                                                                                                                                                                                                                                                                                                                                  V        f�)    �   L   N          O    getA: somador32 port map (a => sum0Out, b => sum0Complement, s => preAOut);�   K   M          a    getSum0Complement: somador32 port map (a => majOut, b => majComplement, s => sum0Complement);�   J   L          I    getE: somador32 port map (a => di, b => majComplement, s => preEOut);�   I   K          a    getMajComplement: somador32 port map (a => sum1Out, b => sum1Complement, s => majComplement);�   H   J          _    getSum1Complement: somador32 port map (a => chOut, b => chComplement, s => sum1Complement);�   G   I          O    getChComplement: somador32 port map (a => hi, b => kpw, s => chComplement);�   &   (   X          component somador32 is5��    &          	          �      	              �    G          	          �      	              �    H          	          �      	              �    I          	          D      	              �    J   
       	          �      	              �    K          	          �      	              �    L   
       	          @	      	              5�_�                            ����                                                                                                                                                                                                                                                                                                                                      W          V       f�     �       Y         entity stepfun is�             �             V   
    port (   @    	ai, bi, ci, di, ei, fi, gi, hi: in bit_vector(31 downto 0);   (        kpw: in bit_vector(31 downto 0);   C        ao, bo, co, do, eo, fo, go, ho: out bit_vector(31 downto 0)   
        );   end stepfun;       %architecture behavioral of stepfun is   #    -- Declaração dos componentes       component ch is           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component maj is           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component sum0 is           port (   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component sum1 is           port (   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component adder32 is           port (   +            a : in bit_vector(31 downto 0);   +            b : in bit_vector(31 downto 0);   +            s : out bit_vector(31 downto 0)   
        );       end component;           -- Sinais           -- Sums complements   1    signal chComplement: bit_vector(31 downto 0);   2    signal majComplement: bit_vector(31 downto 0);   3    signal sum0Complement: bit_vector(31 downto 0);   3    signal sum1Complement: bit_vector(31 downto 0);       "    -- Crytografy funcions outputs   +    signal chOut: bit_vector(31 downto 0);    ,    signal majOut: bit_vector(31 downto 0);    -    signal sum0Out: bit_vector(31 downto 0);    -    signal sum1Out: bit_vector(31 downto 0);            -- Intermediate outputs   ,    signal preAOut: bit_vector(31 downto 0);   ,    signal preEOut: bit_vector(31 downto 0);       begin       -- Saida dos Componentes   +    getCh: ch port map (ei, fi, gi, chOut);   .    getMaj: maj port map (ai, bi, ci, majOut);   )    getSum0: sum0 port map (ai, sum0Out);   )    getSum1: sum1 port map (ei, sum1Out);       M    getChComplement: adder32 port map (a => hi, b => kpw, s => chComplement);   ]    getSum1Complement: adder32 port map (a => chOut, b => chComplement, s => sum1Complement);   _    getMajComplement: adder32 port map (a => sum1Out, b => sum1Complement, s => majComplement);   G    getE: adder32 port map (a => di, b => majComplement, s => preEOut);   _    getSum0Complement: adder32 port map (a => majOut, b => majComplement, s => sum0Complement);   M    getA: adder32 port map (a => sum0Out, b => sum0Complement, s => preAOut);           ao <= preAOut;       bo <= ai;       co <= bi;       do <= ci;       eo <= preEOut;       fo <= ei;       go <= fi;       ho <= gi;   end behavioral;5��           V                      �	              �                                                  �                    W                       
      5�_�                    X        ����                                                                                                                                                                                                                                                                                                                                      Y          V       f�	    �   W   X           5��    W                      
                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                       X           V        f��   	 �                  entity stepfun is�               �             W   
    port (   @    	ai, bi, ci, di, ei, fi, gi, hi: in bit_vector(31 downto 0);   (        kpw: in bit_vector(31 downto 0);   C        ao, bo, co, do, eo, fo, go, ho: out bit_vector(31 downto 0)   
        );   end stepfun;       %architecture behavioral of stepfun is   #    -- Declaração dos componentes       component ch is           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component maj is           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component sum0 is           port (   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component sum1 is           port (   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component somador is           port (   +            A : in bit_vector(31 downto 0);   +            B : in bit_vector(31 downto 0);   +            S : out bit_vector(31 downto 0)   
        );       end component;           -- Sinais           -- Sums complements   1    signal chComplement: bit_vector(31 downto 0);   2    signal majComplement: bit_vector(31 downto 0);   3    signal sum0Complement: bit_vector(31 downto 0);   3    signal sum1Complement: bit_vector(31 downto 0);       "    -- Crytografy funcions outputs   +    signal chOut: bit_vector(31 downto 0);    ,    signal majOut: bit_vector(31 downto 0);    -    signal sum0Out: bit_vector(31 downto 0);    -    signal sum1Out: bit_vector(31 downto 0);            -- Intermediate outputs   ,    signal preAOut: bit_vector(31 downto 0);   ,    signal preEOut: bit_vector(31 downto 0);       begin       -- Saida dos Componentes   +    getCh: ch port map (ei, fi, gi, chOut);   .    getMaj: maj port map (ai, bi, ci, majOut);   )    getSum0: sum0 port map (ai, sum0Out);   )    getSum1: sum1 port map (ei, sum1Out);       M    getChComplement: somador port map (A => hi, B => kpw, S => chComplement);   ]    getSum1Complement: somador port map (A => chOut, B => chComplement, S => sum1Complement);   _    getMajComplement: somador port map (A => sum1Out, B => sum1Complement, S => majComplement);   G    getE: somador port map (A => di, B => majComplement, S => preEOut);   _    getSum0Complement: somador port map (A => majOut, B => majComplement, S => sum0Complement);   M    getA: somador port map (A => sum0Out, B => sum0Complement, S => preAOut);           ao <= preAOut;       bo <= ai;       co <= bi;       do <= ci;       eo <= preEOut;       fo <= ei;       go <= fi;       ho <= gi;   end behavioral;    5��           W                      �	              �                                                  �                    G                      �      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f�     �         H      	component somadorNbits is5��                        4                    5�_�                            ����                                                                                                                                                                                                                                                                                                                               
                 V       f�     �                		generic (   				N		: positive := 32   		);5��                          ?      )               5�_�                           ����                                                                                                                                                                                                                                                                                                                               
                 V       f�"     �         E      +		port (a	 	: in  bit_vector(N-1 downto 0);5��                        G              	       �                         H                    5�_�                           ����                                                                                                                                                                                                                                                                                                                               
                 V       f�#     �         F      4                 a	 	: in  bit_vector(N-1 downto 0);5��                         X                     5�_�                       %    ����                                                                                                                                                                                                                                                                                                                               
                 V       f�(     �         F      3                a	 	: in  bit_vector(N-1 downto 0);5��       %                  m                     5�_�                       %    ����                                                                                                                                                                                                                                                                                                                               
                 V       f�(     �         F      2                a	 	: in  bit_vector(-1 downto 0);5��       %                  m                     5�_�                       %    ����                                                                                                                                                                                                                                                                                                                               
                 V       f�)     �         F      1                a	 	: in  bit_vector(1 downto 0);5��       %                  m                     5�_�                           ����                                                                                                                                                                                                                                                                                                                               
                 V       f�+     �         F      '				b  	: in  bit_vector(N-1 downto 0);5��                         �                     5�_�                            ����                                                                                                                                                                                                                                                                                                                               
                 V       f�,     �         F      &				b  	: in  bit_vector(-1 downto 0);5��                         �                     5�_�      !                      ����                                                                                                                                                                                                                                                                                                                               
                 V       f�-     �         F      %				b  	: in  bit_vector(1 downto 0);5��                         �                     5�_�       "           !          ����                                                                                                                                                                                                                                                                                                                               
                 V       f�/     �                				cin   : in  bit;5��                          �                     5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                               
                 V       f�1     �         E      &				s		: out bit_vector(N-1 downto 0);5��                         �                     �                        �                    5�_�   "   $           #          ����                                                                                                                                                                                                                                                                                                                               
                 V       f�4     �                				cout	: out bit5��                          �                     5�_�   #   %           $      %    ����                                                                                                                                                                                                                                                                                                                               
                 V       f�9     �         D      %				s		: out bit_vector(31 downto 0);5��       $                  �                     5�_�   $               %           ����                                                                                                                                                                                                                                                                                                                               
                 V       f�e   
 �                	component adder32 is   		port (   2                a	 	: in  bit_vector(31 downto 0);   &				b  	: in  bit_vector(31 downto 0);   $				s		: out bit_vector(31 downto 0)   		);   	end component;    5��                          )      �               5�_�                    '        ����                                                                                                                                                                                                                                                                                                                                                             fmw     �   &   (   X          component adder32 is�   G   I          M    getChComplement: adder32 port map (A => hi, B => kpw, S => chComplement);�   H   J          ]    getSum1Complement: adder32 port map (A => chOut, B => chComplement, S => sum1Complement);�   I   K          _    getMajComplement: adder32 port map (A => sum1Out, B => sum1Complement, S => majComplement);�   J   L          G    getE: adder32 port map (A => di, B => majComplement, S => preEOut);�   K   M          _    getSum0Complement: adder32 port map (A => majOut, B => majComplement, S => sum0Complement);�   L   N          M    getA: adder32 port map (A => sum0Out, B => sum0Complement, S => preAOut);5��    &                    �                    �    G                    �                    �    H                    �                    �    I                    D                    �    J   
                 �                    �    K                    �                    �    L   
                 @	                    5��