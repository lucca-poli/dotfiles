Vim�UnDo� ����f�~�
m�LD�oo��-J�^�~ �m   :           !      7       7   7   7    f�C    _�                             ����                                                                                                                                                                                                                                                                                                                                                             fv�     �                   �               5��                   P                      5	      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             fv�     �                  5��                                                  5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             fv�     �   !   #              dut: counter_6bit�                    component counter_6bit�                (architecture Behavioral of counter_tb is�         P      entity counter_tb is end;5��                     
   0              
       �                     
   b              
       �                     
   �              
       �    !   	              
   �             
       5�_�                    "       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   !   #   P          dut: multisteps_6bit5��    !                     �                     5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                             f��     �         P          component multisteps_6bit5��                         �                      5�_�      
           	   	        ����                                                                                                                                                                                                                                                                                                                            	                    V       f��     �         M    �   	   
   M    �      	          C            clk : in bit;                            -- Clock input   A            rst : in bit;                          -- Reset input   U            count : out bit_vector(5 downto 0)       -- 6-bit count output (64 steps)5��                          �       �               �                          �               �       5�_�   	              
   	       ����                                                                                                                                                                                                                                                                                                                            	                           f��     �   	      Q      +        msgi : in bit_vector(511 downto 0);   ,        haso : out bit_vector(255 downto 0);           done : out bit�      
   Q              clk, rst : in bit;5��                         �                      �    	                     �                      �    
                     �                      �                         #                     5�_�   
                        ����                                                                                                                                                                                                                                                                                                                            	                           f�.     �         Q    5��                          �                     �                          �                     5�_�                            ����                                                                                                                                                                                                                                                                                                                            	                           f�/     �         R    5��                          �                     �                          �                     �                          �                     5�_�                            ����                                                                                                                                                                                                                                                                                                                            	                           f�K     �                 5��                          �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         R      =    signal count : bit_vector(5 downto 0);  -- Input stimulus5��                         	                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         R      8    signal  : bit_vector(5 downto 0);  -- Input stimulus5��                         	                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         R      <    signal msgi : bit_vector(5 downto 0);  -- Input stimulus5��                                            5�_�                          ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         S          �         R    5��                          �                     �                                              �                                            5�_�                       *    ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         S      >    signal msgi : bit_vector(511 downto 0);  -- Input stimulus5��       *                  ;                     �       -                  >                     5�_�                       -    ����                                                                                                                                                                                                                                                                                                                            	                           f�     �         S      A    signal msgi : bit_vector(511 downto 0) :=;  -- Input stimulus5��       -                  >                     5�_�                       .    ����                                                                                                                                                                                                                                                                                                                            	                           f�     �         S      B    signal msgi : bit_vector(511 downto 0) := ;  -- Input stimulus5��       .                  ?                     5�_�                       /    ����                                                                                                                                                                                                                                                                                                                            	                           f�     �         S      D    signal msgi : bit_vector(511 downto 0) := ();  -- Input stimulus5��       /                  @                     �       /                 @                    �       /                 @                    �       /                 @                    �       /                 @                    �       /                 @                    5�_�                       ;    ����                                                                                                                                                                                                                                                                                                                            	                           f�     �         S    �         S    5��                          c              R       5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f�     �         T      Q    signal msgi : bit_vector(511 downto 0) := (others => '0');  -- Input stimulus5��                        �                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f�!     �         T      Q    signal msgi : bit_vector(255 downto 0) := (others => '0');  -- Input stimulus5��                        n                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f�,     �         U          �         T    5��                          �                     �                         �                     �                        �                    5�_�                       *    ����                                                                                                                                                                                                                                                                                                                            	                           f�@    �         U      Q    signal haso : bit_vector(255 downto 0) := (others => '0');  -- Input stimulus5��       *                  �                     5�_�                    +       ����                                                                                                                                                                                                                                                                                                                            	                           f�Z     �   *   ,   U                  count => count5��    *                    5                    �    *                     7                     �    *                     6                     �    *                    5                    �    *                    5                    �    *                    5                    5�_�                    +       ����                                                                                                                                                                                                                                                                                                                            	                           f�^     �   ,   .   W                  done�   +   .   V                  haso�   *   -   U                  msgi => count5��    *                    =                    �    *                     >                     �    *                    =                    �    *                    =                    �    *                    =                    �    *                    B                     �    +                     O                     �    +                    O                    �    +                    O                    �    +                    O                    �    +                    S                    �    +                    U                    �    +                     Y                     �    +                     X                     �    +                    W                    �    +                    W                    �    +                    W                    �    +                    \                     �    ,                     i                     �    ,                    j                    �    ,                    i                    �    ,                    i                    �    ,                    i                    �    ,                     s                     �    ,                     r                     �    ,                    q                    �    ,                    q                    �    ,                    q                    5�_�                    4   !    ����                                                                                                                                                                                                                                                                                                                            	                           f�s     �   3   5   W      6        assert false report "BOT count" severity note;5��    3   !                 �                    �    3   !              
   �             
       �    3   !       
          �      
              �    3   !              
   �             
       5�_�                     S   !    ����                                                                                                                                                                                                                                                                                                                            	                           f��     �   R   T   W      6        assert false report "EOT count" severity note;5��    R   !                 _	                    �    R   !              
   _	             
       �    R   !       
          _	      
              �    R   !              
   _	             
       5�_�      !               Q   *    ����                                                                                                                                                                                                                                                                                                                            	                           f��     �   P   Q          H        assert count = "000001" report "Did not proceed" severity error;5��    P                      �      I               5�_�       "           !   O        ����                                                                                                                                                                                                                                                                                                                            	                           f��     �   N   O          &        rst <= '0';  -- Deassert reset5��    N                      �      '               5�_�   !   #           "   L        ����                                                                                                                                                                                                                                                                                                                            	                           f��     �   K   L          $        rst <= '1';  -- Assert reset5��    K                      �      %               5�_�   "   $           #   L        ����                                                                                                                                                                                                                                                                                                                L           	                           f��     �   K   M   T      7        wait for CLOCK_PERIOD;  -- Hold reset for 20 ns   F        assert count = "000000" report "Did not reset" severity error;5��    K   7                (      	              5�_�   #   %           $   L        ����                                                                                                                                                                                                                                                                                                                L           	                           f��     �   K   M   S      v        wait for CLOCK_PERIOD;  -- Hold reset for 20 ns assert count = "000000" report "Did not reset" severity error;   7        wait for CLOCK_PERIOD;  -- Hold reset for 20 ns5��    K   v                g      	              5�_�   $   &           %   7        ����                                                                                                                                                                                                                                                                                                                L           L           7           V        f��     �   6   7          '        assert count = "000001" report    V        "Did not proceed to 1, count is " & integer'image(to_integer(unsigned(count)))           severity error;               wait for CLOCK_PERIOD;   '        assert count = "000010" report    V        "Did not proceed to 2, count is " & integer'image(to_integer(unsigned(count)))           severity error;               wait for CLOCK_PERIOD;   '        assert count = "000011" report    V        "Did not proceed to 3, count is " & integer'image(to_integer(unsigned(count)))           severity error;               wait for CLOCK_PERIOD;   '        assert count = "000100" report    W        "Did not proceed to 4, count is " & integer'image(to_integer(unsigned(count)))            severity error;               wait for CLOCK_PERIOD;       �        wait for CLOCK_PERIOD;  -- Hold reset for 20 ns assert count = "000000" report "Did not reset" severity error; wait for CLOCK_PERIOD;  -- Hold reset for 20 ns5��    6                            �              5�_�   %   '           &   6        ����                                                                                                                                                                                                                                                                                                                            7           7           V        f��     �   6   8   <    �   6   7   <    5��    6                                           5�_�   &   (           '   7       ����                                                                                                                                                                                                                                                                                                                            8           8           V        f��     �   7   9   =    �   7   8   =    5��    7                      2                     5�_�   '   )           (   8       ����                                                                                                                                                                                                                                                                                                                            9           9           V        f��     �   8   :   >    �   8   9   >    5��    8                      Q                     5�_�   (   *           )   9       ����                                                                                                                                                                                                                                                                                                                            :           :           V        f��     �   9   ;   ?    �   9   :   ?    5��    9                      p                     5�_�   )   +           *   :       ����                                                                                                                                                                                                                                                                                                                            ;           ;           V        f��     �   :   <   @    �   :   ;   @    5��    :                      �                     5�_�   *   ,           +   ;       ����                                                                                                                                                                                                                                                                                                                            <           <           V        f��     �   ;   =   A    �   ;   <   A    5��    ;                      �                     5�_�   +   -           ,   <       ����                                                                                                                                                                                                                                                                                                                            =           =           V        f��     �   <   >   B    �   <   =   B    5��    <                      �                     5�_�   ,   .           -   =       ����                                                                                                                                                                                                                                                                                                                            >           >           V        f��     �   =   ?   C    �   =   >   C    5��    =                      �                     5�_�   -   /           .   >       ����                                                                                                                                                                                                                                                                                                                            ?           ?           V        f��     �   >   @   D    �   >   ?   D    5��    >                                           5�_�   .   0           /   ?       ����                                                                                                                                                                                                                                                                                                                            @           @           V        f��     �   ?   A   E    �   ?   @   E    5��    ?                      *                     5�_�   /   1           0   @       ����                                                                                                                                                                                                                                                                                                                            A           A           V        f��     �   @   B   F    �   @   A   F    5��    @                      I                     5�_�   0   2           1   A       ����                                                                                                                                                                                                                                                                                                                            B           B           V        f��     �   A   C   G    �   A   B   G    5��    A                      h                     5�_�   1   3           2   B       ����                                                                                                                                                                                                                                                                                                                            C           C           V        f��     �   B   D   H    �   B   C   H    5��    B                      �                     5�_�   2   4           3   C       ����                                                                                                                                                                                                                                                                                                                            D           D           V        f��    �   C   E   I    �   C   D   I    5��    C                      �                     5�_�   3   6           4   8       ����                                                                                                                                                                                                                                                                                                                            D          8          V       f�*    �   7   8                  wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;           wait for CLOCK_PERIOD;5��    7                      2      �              5�_�   4   7   5       6   6        ����                                                                                                                                                                                                                                                                                                                            8          8          V       f�:    �   5   6                  wait for CLOCK_PERIOD;5��    5                      �                     5�_�   6               7   6        ����                                                                                                                                                                                                                                                                                                                            7          7          V       f�B    �   5   6                  wait for CLOCK_PERIOD;    5��    5                      �                      5�_�   4           6   5   6        ����                                                                                                                                                                                                                                                                                                                            6          6          V       f�8     �   5   8        5��    5                      �      >               5�_�                           ����                                                                                                                                                                                                                                                                                                                            	                           f��     �         R       5��                          =                     �                          =                     5�_�                          ����                                                                                                                                                                                                                                                                                                                                                             fv�     �         P      entity mul_tb is end;5��                        0                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             fv�     �               5��                                                  5�_�                             ����                                                                                                                                                                                                                                                                                                                                                             fv�     �               5��                                                  5��