Vim�UnDo� �#�DuM�P�s6���ta(t��D���OC�   \           wait;   Z                          f(�    _�                     Z       ����                                                                                                                                                                                                                                                                                                                                                             f(�     �   Y   [   \              wait for 1ms;5��    Y                     �
                     5�_�                     Z       ����                                                                                                                                                                                                                                                                                                                                                             f(�    �   Y   [   \              wait for 1 ms;5��    Y                     �
                     5��