Vim�UnDo� B�^+[Y���V��v6���@�2�XrhD��m8<   �   c            " Computed Q=" & to_hstring(unsigned(ho)) & ", Expected Q=" & to_hstring(unsigned(Hov))   }         �       �   �   �    fٱ   
 _�                             ����                                                                                                                                                                                                                                                                                                                                                             e��$     �                >        file tb_file : text open read_mode is "cases/maj.dat";�                    dut: maj�      
              component maj�                architecture dut of maj_tb is�         G      entity maj_tb is end;5��                        D                     �                        i                     �                        �                     �       	                 �                    �       5                 �                    5�_�                    1        ����                                                                                                                                                                                                                                                                                                                            ,          .          V       e��?     �   1   5   G    �   1   2   G    5��    1                      �              V       5�_�                    4       ����                                                                                                                                                                                                                                                                                                                            ,          .          V       e��@     �   4   8   J    �   4   5   J    5��    4                      F              V       5�_�                    7       ����                                                                                                                                                                                                                                                                                                                            ,          .          V       e��B     �   7   ;   M    �   7   8   M    5��    7                      �              V       5�_�                    :       ����                                                                                                                                                                                                                                                                                                                            ,          .          V       e��C     �   :   >   P    �   :   ;   P    5��    :                      �              V       5�_�      
              =       ����                                                                                                                                                                                                                                                                                                                            ,          .          V       e��D     �   =   A   S    �   =   >   S    5��    =                      H              V       5�_�                
          ����                                                                                                                                                                                                                                                                                                                            ,          .          V       e��h     �         V      6        port map (x => x, y => y, z => z, q => saida);5��                                      	       �                                             5�_�   
                        ����                                                                                                                                                                                                                                                                                                                            -          /          V       e��k     �         W      .                  y => y, z => z, q => saida);5��                        /                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            .          0          V       e��m     �         X      &                  z => z, q => saida);5��                        J                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          1          V       e��t     �         Y      -    signal x, y, z : bit_vector(31 downto 0);5��                        z                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          1          V       e��v     �         Y      .    signal ai, y, z : bit_vector(31 downto 0);5��                        ~                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          1          V       e��y     �         Y      /    signal ai, bi, z : bit_vector(31 downto 0);5��                        �                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          1          V       e��}     �         Y      +    signal saida : bit_vector(31 downto 0);5��                        �                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          1          V       e�ڎ     �         Y      0    signal ai, bi, ci : bit_vector(31 downto 0);5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          1          V       e�ڝ     �         Y              port map (x => x, 5��                        A                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          1          V       e�ڟ     �         Y              port map (ai => x, 5��                        G                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          1          V       e�ڢ     �         Y                        y => y, 5��                        ^                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          1          V       e�ڤ     �         Y                        bi => y, 5��                        d                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          1          V       e�ڧ     �         Y                        z => z, 5��                        {                    �                        {                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          1          V       e�ک     �         Y                        ci => z, 5��                        �                    �                         �                     �                        �                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          1          V       e�ڳ     �         Y                        bi => ci, 5��                        d                    5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          1          V       e�ڵ     �         Y    �         Y    5��                          �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            0          2          V       e�ڶ     �         Z    �         Z    5��                          �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            1          3          V       e�ڷ     �         [    �         [    5��                          �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            2          4          V       e�ڸ     �         \    �         \    5��                          �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            3          5          V       e�ڸ     �          ]    �         ]    5��                          �                     5�_�                            ����                                                                                                                                                                                                                                                                                                                            4          6          V       e��     �         ^                        ci => ci, 5�5�_�      !                     ����                                                                                                                                                                                                                                                                                                                            4          6          V       e��5     �         ^                        ci => ci, 5�5�_�       "           !           ����                                                                                                                                                                                                                                                                                                                                                  V        e�ݱ     �         ^                        ci => ci, 5��                        �                    �                        �                    5�_�   !   #           "           ����                                                                                                                                                                                                                                                                                                                                                V       e���     �         ^                        ci => ci, 5��                        �                    �                        �                    5�_�   "   $           #           ����                                                                                                                                                                                                                                                                                                                                                V       e���     �         ^                        ci => ci, 5��                        �                    �                        �                    5�_�   #   %           $           ����                                                                                                                                                                                                                                                                                                                                                V       e���     �         ^                        di => di, 5��                        �                    �                        �                    5�_�   $   &           %           ����                                                                                                                                                                                                                                                                                                                                                V       e���     �         ^                        di => di, 5��                        �                    �                        �                    �                        �                    �                        �                    5�_�   %   '           &           ����                                                                                                                                                                                                                                                                                                                                                V       e���     �         ^                        ci => ci, 5��                        �                    �                        �                    �                        �                    �                        �                    �                        �                    �                        �                    5�_�   &   (           '           ����                                                                                                                                                                                                                                                                                                                                                V       e���     �          ^                        ci => ci, 5��                                            �                                            �                                            �                                            �                                            �                                            �                                            �                                            5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                V       e��      �                                  gi => gi, 5��                          �                     5�_�   (   *           )          ����                                                                                                                                                                                                                                                                                                                                                V       e��     �         ]    �         ]    5��                          �                     5�_�   )   +           *           ����                                                                                                                                                                                                                                                                                                                                                V       e��     �          ^                        fi => fi, 5��                                            �                                            �                                            �                                            5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                                V       e��     �      !   ^    �          ^    5��                                               5�_�   +   -           ,           ����                                                                                                                                                                                                                                                                                                                                                V       e��     �      !   _                        hi => hi, 5��                        )                    5�_�   ,   .           -           ����                                                                                                                                                                                                                                                                                                                                                V       e��     �      !   _                        kpw => hi, 5��                        0                    5�_�   -   3           .           ����                                                                                                                                                                                                                                                                                                                                                V       e��     �       "   _    �       !   _    5��                           6                     5�_�   .   4   /       3   !       ����                                                                                                                                                                                                                                                                                                                                                V       e��     �       "   `                        hi => hi, 5��                          I                     �                         H                    5�_�   3   5           4   !       ����                                                                                                                                                                                                                                                                                                                                                V       e��     �       "   `                        ai => hi, 5��                         N                    5�_�   4   6           5   !       ����                                                                                                                                                                                                                                                                                                                                                V       e��!     �       "   `                        ai => ao, 5��                         I                    5�_�   5   7           6   !       ����                                                                                                                                                                                                                                                                                                                                                V       e��"     �       "   `                        a0 => ao, 5��                         I                    5�_�   6   8           7   !       ����                                                                                                                                                                                                                                                                                                                                                V       e��#     �   !   #   `    �   !   "   `    5��    !                      S                     5�_�   7   9           8   "       ����                                                                                                                                                                                                                                                                                                                                                V       e��$     �   "   $   a    �   "   #   a    5��    "                      p                     5�_�   8   :           9   #       ����                                                                                                                                                                                                                                                                                                                                                V       e��%     �   #   %   b    �   #   $   b    5��    #                      �                     5�_�   9   ;           :   $       ����                                                                                                                                                                                                                                                                                                                                                V       e��&     �   $   &   c    �   $   %   c    5��    $                      �                     5�_�   :   <           ;   %       ����                                                                                                                                                                                                                                                                                                                                                V       e��&     �   %   '   d    �   %   &   d    5��    %                      �                     5�_�   ;   =           <   &       ����                                                                                                                                                                                                                                                                                                                                                V       e��&     �   &   (   e    �   &   '   e    5��    &                      �                     5�_�   <   >           =   '       ����                                                                                                                                                                                                                                                                                                                                                V       e��'     �   '   )   f    �   '   (   f    5��    '                                           5�_�   =   ?           >   (       ����                                                                                                                                                                                                                                                                                                                                                V       e��'     �   (   *   g    �   (   )   g    5��    (                                           5�_�   >   @           ?   )       ����                                                                                                                                                                                                                                                                                                                                                V       e��*     �   (   )                            ao => ao, 5��    (                                           5�_�   ?   A           @   )       ����                                                                                                                                                                                                                                                                                                                                                V       e��0     �   '   )   g                        ao => ao,    );�   (   *   g                        q => saida);5��    (                                           �    '                                          �    '                                          �    '                                          5�_�   @   B           A   "        ����                                                                                                                                                                                                                                                                                                                            "          "          V       e��7     �   !   #   f                        ao => ao, 5��    !                    e                    �    !                    k                    5�_�   A   C           B   #        ����                                                                                                                                                                                                                                                                                                                            #          #          V       e��:     �   "   $   f                        ao => ao, 5��    "                    �                    �    "                    �                    �    "                    �                    �    "                    �                    5�_�   B   D           C   $        ����                                                                                                                                                                                                                                                                                                                            $          $          V       e��<     �   #   %   f                        ao => ao, 5��    #                    �                    �    #                    �                    �    #                    �                    �    #                    �                    �    #                    �                    �    #                    �                    5�_�   C   E           D   %        ����                                                                                                                                                                                                                                                                                                                            %          %          V       e��>     �   $   &   f                        ao => ao, 5��    $                    �                    �    $                    �                    �    $                    �                    �    $                    �                    �    $                    �                    �    $                    �                    �    $                    �                    �    $                    �                    5�_�   D   F           E   &        ����                                                                                                                                                                                                                                                                                                                            &          &          V       e��@     �   %   '   f                        ao => ao, 5��    %                    �                    �    %                    �                    �    %                    �                    �    %                    �                    �    %                    �                    �    %                    �                    �    %                    �                    �    %                    �                    �    %                    �                    �    %                    �                    5�_�   E   G           F   '        ����                                                                                                                                                                                                                                                                                                                            '          '          V       e��C     �   &   (   f                        ao => ao, 5��    &                    �                    �    &                    �                    �    &                    �                    �    &                    �                    �    &                    �                    �    &                    �                    �    &                    �                    �    &                    �                    �    &                    �                    �    &                    �                    �    &                    �                    �    &                    �                    5�_�   F   H           G   (        ����                                                                                                                                                                                                                                                                                                                            (          (          V       e��E    �   '   )   f                        ao => ao);5��    '                                        �    '                                        �    '                                        �    '                                        �    '                                        �    '                                        �    '                                        �    '                                        �    '                                        �    '                                        �    '                                        �    '                                        �    '                                        �    '                                        5�_�   G   I           H          ����                                                                                                                                                                                                                                                                                                                                                V       e�ބ     �   
      d    �         d    �   
             0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)5��    
                      �       \               �    
                      �               �       5�_�   H   K           I          ����                                                                                                                                                                                                                                                                                                                                                       e�ވ     �         g      (        kpw: in bit_vector(31 downto 0);   C        ao, bo, co, do, eo, fo, go, ho: out bit_vector(31 downto 0)�   
      g      @    	ai, bi, ci, di, ei, fi, gi, hi: in bit_vector(31 downto 0);5��    
                     �                      �                                               �                         M                     5�_�   I   L   J       K   0       ����                                                                                                                                                                                                                                                                                                                                                       e�ޘ     �   /   1   g      :        variable Xv, Yv, Zv, res: bit_vector(31 downto 0);5��    /                    >                    5�_�   K   M           L   0       ����                                                                                                                                                                                                                                                                                                                                                       e�ޚ     �   /   1   g      :        variable Av, Yv, Zv, res: bit_vector(31 downto 0);5��    /                     ?                     5�_�   L   N           M   0       ����                                                                                                                                                                                                                                                                                                                                                       e�ި     �   /   1   g      ;        variable Aiv, Yv, Zv, res: bit_vector(31 downto 0);5��    /                    C                    5�_�   M   O           N   0       ����                                                                                                                                                                                                                                                                                                                                                       e�ޫ     �   /   1   g      <        variable Aiv, Biv, Zv, res: bit_vector(31 downto 0);5��    /                    H                    5�_�   N   P           O   0        ����                                                                                                                                                                                                                                                                                                                                                       e�ޮ     �   /   1   g      =        variable Aiv, Biv, Civ, res: bit_vector(31 downto 0);5��    /                     M                    5�_�   O   Q           P   0   #    ����                                                                                                                                                                                                                                                                                                                                                       e�޳     �   /   1   g      =        variable Aiv, Biv, Civ, Div: bit_vector(31 downto 0);5��    /   #                  P                     �    /   6                 c                    �    /   7                 d                    5�_�   P   R           Q   0   <    ����                                                                                                                                                                                                                                                                                                                                                       e���     �   0   2   g    �   0   1   g    5��    0                      �              X       5�_�   Q   S           R   1        ����                                                                                                                                                                                                                                                                                                                            1          1          V       e���     �   0   2   h      W        variable Aiv, Biv, Civ, Div, Eiv, Fiv, Giv, Hiv, KpwV: bit_vector(31 downto 0);5��    0                    �                    �    0                    �                    �    0                    �                    �    0                    �                    �    0   !                 �                    �    0   &                 �                    �    0   +                 �                    �    0   0                 �                    �    0   5                 �                    �    0   @                 �                    5�_�   R   T           S   1       ����                                                                                                                                                                                                                                                                                                                            1          1          V       e���     �   0   2   h      W        varoable Aov, Bov, Cov, Dov, Eov, Fov, Gov, Hov, KpwV: bot_vector(31 downto 0);5��    0                    �                    5�_�   S   U           T   1   9    ����                                                                                                                                                                                                                                                                                                                            1          1          V       e���     �   0   2   h      W        variable Aov, Bov, Cov, Dov, Eov, Fov, Gov, Hov, KpwV: bot_vector(31 downto 0);5��    0   9                  �                     5�_�   T   V           U   1   7    ����                                                                                                                                                                                                                                                                                                                            1          1          V       e���     �   0   2   h      S        variable Aov, Bov, Cov, Dov, Eov, Fov, Gov, Hov, : bot_vector(31 downto 0);5��    0   7                  �                     5�_�   U   W           V   1   7    ����                                                                                                                                                                                                                                                                                                                            1          1          V       e���     �   0   2   h      R        variable Aov, Bov, Cov, Dov, Eov, Fov, Gov, Hov : bot_vector(31 downto 0);5��    0   7                  �                     5�_�   V   X           W   1   :    ����                                                                                                                                                                                                                                                                                                                            1          1          V       e���     �   0   2   h      Q        variable Aov, Bov, Cov, Dov, Eov, Fov, Gov, Hov: bot_vector(31 downto 0);5��    0   :                 �                    5�_�   W   Y           X   <       ����                                                                                                                                                                                                                                                                                                                            1          1          V       e���     �   ;   =   h                  x <= Xv;5��    ;                    �                    5�_�   X   Z           Y   <       ����                                                                                                                                                                                                                                                                                                                            1          1          V       e���     �   ;   =   h                  A <= Xv;5��    ;                    �                    5�_�   Y   [           Z   ;       ����                                                                                                                                                                                                                                                                                                                            1          1          V       e���     �   :   <   h                  read(tb_line, Xv);5��    :                    �                    5�_�   Z   \           [   <       ����                                                                                                                                                                                                                                                                                                                            1          1          V       e���     �   ;   =   h                  ai <= Xv;5��    ;                    �                    5�_�   [   ]           \   >       ����                                                                                                                                                                                                                                                                                                                            1          1          V       e���     �   =   ?   h                  read(tb_line, Yv);5��    =                                        5�_�   \   ^           ]   ?       ����                                                                                                                                                                                                                                                                                                                            1          1          V       e���     �   >   @   h                  y <= Yv;5��    >                    2                    5�_�   ]   _           ^   ?       ����                                                                                                                                                                                                                                                                                                                            1          1          V       e��     �   >   @   h                  y <= Biv;5��    >                    -                    5�_�   ^   `           _   B       ����                                                                                                                                                                                                                                                                                                                            1          1          V       e��     �   A   C   h                  z <= Zv;5��    A                    �                    5�_�   _   a           `   E       ����                                                                                                                                                                                                                                                                                                                            1          1          V       e��     �   D   F   h                  y <= Yv;5��    D                    �                    5�_�   `   b           a   H       ����                                                                                                                                                                                                                                                                                                                            1          1          V       e��	     �   G   I   h                  y <= Yv;5��    G                    3                    5�_�   a   c           b   K       ����                                                                                                                                                                                                                                                                                                                            1          1          V       e��     �   J   L   h                  y <= Yv;5��    J                    �                    �    J                    �                    5�_�   b   d           c   N       ����                                                                                                                                                                                                                                                                                                                            1          1          V       e��     �   M   O   h                  y <= Yv;5��    M                    �                    5�_�   c   e           d   Q       ����                                                                                                                                                                                                                                                                                                                            1          1          V       e��     �   P   R   h                  y <= Yv;5��    P                    8	                    5�_�   d   f           e   R        ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��     �   R   V   h    �   R   S   h    5��    R                      d	              W       5�_�   e   g           f   T       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��     �   S   U   k                  hi <= Yv;5��    S                     �	                     �    S                    �	                    5�_�   f   h           g   A       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��'     �   @   B   k                  read(tb_line, Zv);5��    @                    t                    5�_�   g   i           h   B       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��*     �   A   C   k                  ci <= Zv;5��    A                    �                    5�_�   h   j           i   D       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��-     �   C   E   k                  read(tb_line, Yv);5��    C                    �                    5�_�   i   k           j   E       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��/     �   D   F   k                  di <= Yv;5��    D                    �                    5�_�   j   l           k   E       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��0     �   D   F   k                  di <= DIv;5��    D                    �                    5�_�   k   m           l   G       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��3     �   F   H   k                  read(tb_line, Yv);5��    F                    &                    5�_�   l   n           m   H       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��5     �   G   I   k                  ei <= Yv;5��    G                    >                    �    G                    >                    5�_�   m   o           n   J       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��9     �   I   K   k                  read(tb_line, Yv);5��    I                                        5�_�   n   p           o   K       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��<     �   J   L   k                  fi <= Yv;5��    J                    �                    5�_�   o   q           p   M       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��?     �   L   N   k                  read(tb_line, Yv);5��    L                    �                    5�_�   p   r           q   N       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��B     �   M   O   k                  gi <= Yv;5��    M                    �                    5�_�   q   s           r   P       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��D     �   O   Q   k                  read(tb_line, Yv);5��    O                    1	                    5�_�   r   t           s   Q       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��G     �   P   R   k                  hi <= Yv;5��    P                    I	                    5�_�   s   u           t   S       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��K     �   R   T   k                  read(tb_line, Yv);5��    R                    �	                    5�_�   t   v           u   T       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��W     �   S   U   k                  kpw <= Yv;5��    S                    �	                    5�_�   u   w           v   V       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��m     �   V   X   k    �   V   W   k    5��    V                      �	              "       5�_�   v   x           w   V       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e��o     �   U   W   l                  read(tb_line, res);5��    U                    �	                    �    U                     �	                     �    U                     �	                     5�_�   w   y           x   V       ����                                                                                                                                                                                                                                                                                                                            P          R          V       e�߃     �   U   W   l                  read(tb_line, );5��    U                     �	                     5�_�   x   z           y   W        ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�߈     �   W   Z   l    �   W   X   l    5��    W                      
              B       5�_�   y   |           z   Y       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߊ     �   Y   \   n    �   Y   Z   n    5��    Y                      P
              B       5�_�   z   }   {       |   [        ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߍ     �   [   ^   p    �   [   \   p    5��    [                      �
              B       5�_�   |   ~           }   ]       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߎ     �   ]   `   r    �   ]   ^   r    5��    ]                      �
              B       5�_�   }              ~   _       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߏ     �   _   b   t    �   _   `   t    5��    _                                    B       5�_�   ~   �              a       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߏ     �   a   d   v    �   a   b   v    5��    a                      X              B       5�_�      �           �   c       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߐ     �   c   f   x    �   c   d   x    5��    c                      �              B       5�_�   �   �           �   X       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߖ     �   W   Y   z                  read(tb_line, Aov);5��    W                    (
                    5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߘ     �   Y   [   z                  read(tb_line, Aov);5��    Y                    j
                    5�_�   �   �           �   \       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߙ     �   [   ]   z                  read(tb_line, Aov);5��    [                    �
                    5�_�   �   �           �   ^       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߛ     �   ]   _   z                  read(tb_line, Aov);5��    ]                    �
                    5�_�   �   �           �   `       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߝ     �   _   a   z                  read(tb_line, Aov);5��    _                    0                    5�_�   �   �           �   b       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߞ     �   a   c   z                  read(tb_line, Aov);5��    a                    r                    5�_�   �   �           �   d       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߠ     �   c   e   z                  read(tb_line, Aov);5��    c                    �                    5�_�   �   �           �   i       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߵ     �   h   k   z      %            assert saida = res report5��    h                                         5�_�   �   �           �   j       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�߸     �   i   l   {                  saida = res report5��    i                    %                     5�_�   �   �           �   j       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߺ     �   i   k   |                  saida = res 5��    i                                        5�_�   �   �           �   j       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�߾     �   i   k   |                  Aov = res 5��    i                                        5�_�   �   �           �   e       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   d   e          !            read(tb_line, space);5��    d                      �      "               5�_�   �   �           �   i       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   h   j   {                  Aov = ao 5��    h                     �                     5�_�   �   �           �   i       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   h   j   {                  (Aov = ao 5��    h                     �                    5�_�   �   �           �   i       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   h   j   {                  (Aov = ao )5��    h                                           5�_�   �   �           �   i       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   h   j   {                  (Aov = ao)5��    h                                          5�_�   �   �           �   i       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   i   k   {    �   i   j   {    5��    i                                           5�_�   �   �           �   j       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   j   l   |    �   j   k   |    5��    j                      !                     5�_�   �   �           �   k       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   k   m   }    �   k   l   }    5��    k                      <                     5�_�   �   �           �   l       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   l   n   ~    �   l   m   ~    5��    l                      W                     5�_�   �   �           �   m       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   m   o       �   m   n       5��    m                      r                     5�_�   �   �           �   n       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   n   p   �    �   n   o   �    5��    n                      �                     5�_�   �   �           �   o       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   o   q   �    �   o   p   �    5��    o                      �                     5�_�   �   �           �   p       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   o   q   �                  (Aov = ao) and5��    o                     �                     5�_�   �   �           �   j       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   i   k   �                  (Aov = ao) and5��    i                                        5�_�   �   �           �   j       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   i   k   �                  (Bov = ao) and5��    i                                        5�_�   �   �           �   k       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   j   l   �                  (Aov = ao) and5��    j                    4                    5�_�   �   �           �   k       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   j   l   �                  (Aov = jo) and5��    j                    4                    5�_�   �   �           �   l       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   k   m   �                  (Aov = ao) and5��    k                    O                    5�_�   �   �           �   m       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   l   n   �                  (Aov = ao) and5��    l                    j                    5�_�   �   �           �   n       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   m   o   �                  (Aov = ao) and5��    m                    �                    5�_�   �   �           �   o       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   n   p   �                  (Aov = ao) and5��    n                    �                    5�_�   �   �           �   p       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   o   q   �                  (Aov = ao)5��    o                    �                    5�_�   �   �           �   k       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   j   l   �                  (Aov = co) and5��    j                    .                    5�_�   �   �           �   l       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   k   m   �                  (Aov = do) and5��    k                    I                    5�_�   �   �           �   m       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   l   n   �                  (Aov = eo) and5��    l                    d                    5�_�   �   �           �   n       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   m   o   �                  (Aov = fo) and5��    m                                        5�_�   �   �           �   o       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   n   p   �                  (Aov = go) and5��    n                    �                    5�_�   �   �           �   p       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e���     �   o   q   �                  (Aov = ho)5��    o                    �                    5�_�   �   �   �       �   u       ����                                                                                                                                                                                                                                                                                                                            s          u          V       e��     �   r   v   �      =            " X=" & integer'image(to_integer(signed(x))) &LF&   =            " Y=" & integer'image(to_integer(signed(y))) &LF&   =            " Z=" & integer'image(to_integer(signed(z))) &LF&5��    r                     �      �       �       5�_�   �   �           �   v   =    ����                                                                                                                                                                                                                                                                                                                            s          u          V       e��     �   u   w   �      J            " Computed Q=" & integer'image(to_integer(signed(saida))) &LF&5��    u   =                 �                    5�_�   �   �           �   v   @    ����                                                                                                                                                                                                                                                                                                                            s          u          V       e��D     �   u   w   �      H            " Computed Q=" & integer'image(to_integer(signed(Aov))) &LF&5��    u   =                 �                    5�_�   �   �           �   w   =    ����                                                                                                                                                                                                                                                                                                                            s          u          V       e��F    �   v   x   �      C            " Expected Q=" & integer'image(to_integer(signed(res)))5��    v   =                 ;                    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            s          u          V       e���    �   ,   .          ?        file tb_file : text open read_mode is "cases/exp3.dat";�                    dut: exp3�      
              component exp3�                architecture dut of exp3_tb is�         �      entity exp3_tb is end;5��                        D                     �                        l                     �                        �                     �       	                 �                    �    ,   5                 �                    5�_�   �   �   �       �      	    ����                                                                                                                                                                                                                                                                                                                            s          u          V       e���    �               �   library ieee;   use std.textio.all;   use ieee.numeric_bit.ALL;       entity stepfun_tb is end;       !architecture dut of stepfun_tb is   <    -- Component declaration for the DUT (Design Under Test)       component stepfun           port (   D    	    ai, bi, ci, di, ei, fi, gi, hi: in bit_vector(31 downto 0);   ,            kpw: in bit_vector(31 downto 0);   G            ao, bo, co, do, eo, fo, go, ho: out bit_vector(31 downto 0)   
        );       end component;            -- Signals for the testbench   I    signal ai, bi, ci, di, ei, fi, gi, hi, kpw : bit_vector(31 downto 0);   D    signal ao, bo, co, do, eo, fo, go, ho : bit_vector(31 downto 0);       begin           -- Instantiate the DUT       dut: stepfun           port map (ai => ai,                      bi => bi,                      ci => ci,                      di => di,                      ei => ei,                      fi => fi,                      gi => gi,                      hi => hi,                      kpw => kpw,                      ao => ao,                      bo => bo,                      co => co,                      do => do,                      eo => eo,                      fo => fo,                      go => go,                      ho => ho);           -- Stimulus process       stim: process is   B        file tb_file : text open read_mode is "cases/stepfun.dat";           variable tb_line: line;   "        variable space: character;   W        variable Aiv, Biv, Civ, Div, Eiv, Fiv, Giv, Hiv, KpwV: bit_vector(31 downto 0);   Q        variable Aov, Bov, Cov, Dov, Eov, Fov, Gov, Hov: bit_vector(31 downto 0);       	    begin           -- Início do teste   <        assert false report "BOT ch function" severity note;       '        while not endfile(tb_file) loop               -- read inputs   '            readline(tb_file, tb_line);                   read(tb_line, Aiv);               ai <= Aiv;   !            read(tb_line, space);               read(tb_line, Biv);               bi <= Biv;   !            read(tb_line, space);               read(tb_line, Civ);               ci <= Civ;   !            read(tb_line, space);               read(tb_line, Div);               di <= Div;   !            read(tb_line, space);               read(tb_line, Eiv);               ei <= Eiv;   !            read(tb_line, space);               read(tb_line, Fiv);               fi <= Fiv;   !            read(tb_line, space);               read(tb_line, Giv);               gi <= Giv;   !            read(tb_line, space);               read(tb_line, Hiv);               hi <= Hiv;   !            read(tb_line, space);                read(tb_line, Kpwv);               kpw <= Kpwv;   !            read(tb_line, space);               read(tb_line, Aov);   !            read(tb_line, space);               read(tb_line, Bov);   !            read(tb_line, space);               read(tb_line, Cov);   !            read(tb_line, space);               read(tb_line, Dov);   !            read(tb_line, space);               read(tb_line, Eov);   !            read(tb_line, space);               read(tb_line, Fov);   !            read(tb_line, space);               read(tb_line, Gov);   !            read(tb_line, space);               read(tb_line, Hov);                   wait for 1 ns;                   assert                (Aov = ao) and               (Bov = bo) and               (Cov = co) and               (Dov = do) and               (Eov = eo) and               (Fov = fo) and               (Gov = go) and               (Hov = ho)               report                "Output failed" &LF&   @            -- " X=" & integer'image(to_integer(signed(x))) &LF&   @            -- " Y=" & integer'image(to_integer(signed(y))) &LF&   @            -- " Z=" & integer'image(to_integer(signed(z))) &LF&   G            " Computed Q=" & integer'image(to_integer(signed(ao))) &LF&   C            " Expected Q=" & integer'image(to_integer(signed(Aov)))               severity error;               end loop;               -- Fim do teste   <        assert false report "EOT ch function" severity note;       A        wait; -- Wait indefinitely to keep the simulation running       end process;   end dut;    5�5�_�   �   �   �       �   v   6    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   u   w   �      G            " Computed Q=" & integer'image(to_integer(signed(ao))) &LF&5��    u   6                 �                    5�_�   �   �           �   w   6    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   v   x   �      C            " Expected Q=" & integer'image(to_integer(signed(Aov)))5��    v   6                 E                    5�_�   �   �           �   v   .    ����                                                                                                                                                                                                                                                                                                                            w   .       v   4          4    f��     �   u   w   �      B            " Computed Q=" & integer'image(to_(unsigned(ao))) &LF&�   u   x   �      I            " Computed Q=" & integer'image(to_integer(unsigned(ao))) &LF&   E            " Expected Q=" & integer'image(to_integer(unsigned(Aov)))5��    u   .                  �                     �    v   .                  6                     �    u   .                  �                     �    v   .                  =                     5�_�   �   �           �   v       ����                                                                                                                                                                                                                                                                                                                            v          w   *          *    f��     �   u   x   �      I            " Computed Q=" & integer'image(to_hstring(unsigned(ao))) &LF&   E            " Expected Q=" & integer'image(to_hstring(unsigned(Aov)))5��    u                     �                     �    v                                          5�_�   �   �           �   v   4    ����                                                                                                                                                                                                                                                                                                                            v          w   *          *    f��     �   u   w   �      ;            " Computed Q=" & to_hstring(unsigned(ao))) &LF&5��    u   4                  �                     5�_�   �   �           �   w   4    ����                                                                                                                                                                                                                                                                                                                            v          w   *          *    f��    �   v   x   �      7            " Expected Q=" & to_hstring(unsigned(Aov)))5��    v   4                  4                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            v          w   *          *    f�+     �                use ieee.numeric_bit.ALL;5��                          "                      5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            u          v   *          *    f�,    �         �    �         �    5��                                                5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            v          w   *          *    f�K    �         �      use ieee.numeric_bit.ALL;5��                                                5�_�   �   �           �   v   6    ����                                                                                                                                                                                                                                                                                                                            w          w   5       v   5    f�3     �   u   w   �      :            " Computed Q=" & to_hstring(unsigned(ao)) &LF&5��    u   6                  �                     5�_�   �   �           �   v   5    ����                                                                                                                                                                                                                                                                                                                            w          w   5       v   5    f�4     �   u   w   �      ;            " Computed Q=" & to_hstring(unsigned(ao))  &LF&�   v   w   �    5��    u   6               *   �              *       5�_�   �   �           �   v   6    ����                                                                                                                                                                                                                                                                                                                            w          w   5       v   5    f�8     �   u   w   �      e            " Computed Q=" & to_hstring(unsigned(ao)) " Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    u   6                  �                     5�_�   �   �           �   v   9    ����                                                                                                                                                                                                                                                                                                                            w          w   5       v   5    f�:     �   u   w   �      g            " Computed Q=" & to_hstring(unsigned(ao)) & " Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    u   9                                       �    u   :                                       5�_�   �   �           �   w   5    ����                                                                                                                                                                                                                                                                                                                            w          w   5       v   5    f�?     �   v   w          6            " Expected Q=" & to_hstring(unsigned(Aov))5��    v                      2      7               5�_�   �   �   �       �   v       ����                                                                                                                                                                                                                                                                                                                            w          w   5       v   5    f�G     �   v   ~   �    �   v   w   �    5��    v                      2              �      5�_�   �   �           �   w   1    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�N     �   v   x   �      h            " Computed Q=" & to_hstring(unsigned(ao)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    v   1                 c                    5�_�   �   �           �   x   1    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�O     �   w   y   �      h            " Computed Q=" & to_hstring(unsigned(ao)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    w   1                 �                    5�_�   �   �           �   y   1    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�P     �   x   z   �      h            " Computed Q=" & to_hstring(unsigned(ao)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    x   1                 5                    5�_�   �   �           �   y   1    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�Q     �   x   z   �      h            " Computed Q=" & to_hstring(unsigned(fo)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    x   1                 5                    5�_�   �   �           �   z   1    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�S     �   y   {   �      h            " Computed Q=" & to_hstring(unsigned(ao)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    y   1                 �                    5�_�   �   �           �   {   1    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�T     �   z   |   �      h            " Computed Q=" & to_hstring(unsigned(ao)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    z   1                                     5�_�   �   �           �   |   1    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�U     �   {   }   �      h            " Computed Q=" & to_hstring(unsigned(ao)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    {   1                 p                    5�_�   �   �           �   |   1    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�U     �   {   }   �      h            " Computed Q=" & to_hstring(unsigned(go)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    {   1                 p                    5�_�   �   �           �   |   1    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�V     �   {   }   �      h            " Computed Q=" & to_hstring(unsigned(jo)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    {   1                 p                    5�_�   �   �           �   }   1    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�W     �   |   ~   �      h            " Computed Q=" & to_hstring(unsigned(ao)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    |   1                 �                    5�_�   �   �           �   w   ^    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�_     �   v   x   �      h            " Computed Q=" & to_hstring(unsigned(bo)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    v   ^                 �                    5�_�   �   �           �   x   ^    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�`     �   w   y   �      h            " Computed Q=" & to_hstring(unsigned(co)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    w   ^                 �                    5�_�   �   �           �   y   ^    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�a     �   x   z   �      h            " Computed Q=" & to_hstring(unsigned(do)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    x   ^                 b                    5�_�   �   �           �   z   ^    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�b     �   y   {   �      h            " Computed Q=" & to_hstring(unsigned(eo)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    y   ^                 �                    5�_�   �   �           �   {   ^    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�d     �   z   |   �      h            " Computed Q=" & to_hstring(unsigned(fo)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    z   ^                 4                    5�_�   �   �           �   |   ^    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�e     �   {   }   �      h            " Computed Q=" & to_hstring(unsigned(go)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    {   ^                 �                    5�_�   �   �           �   }   ^    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�g     �   |   ~   �      h            " Computed Q=" & to_hstring(unsigned(ho)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    |   ^                                     5�_�   �   �           �   }   d    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�j     �   |   ~   �      h            " Computed Q=" & to_hstring(unsigned(ho)) & ", Expected Q=" & to_hstring(unsigned(Hov)) &LF&5��    |   d                                       5�_�   �   �           �   }   d    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�k     �   |   ~   �      g            " Computed Q=" & to_hstring(unsigned(ho)) & ", Expected Q=" & to_hstring(unsigned(Hov)) LF&5��    |   d                                       5�_�   �   �           �   }   d    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�k     �   |   ~   �      e            " Computed Q=" & to_hstring(unsigned(ho)) & ", Expected Q=" & to_hstring(unsigned(Hov)) &5��    |   d                                       5�_�   �   �           �   }   c    ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f�l   	 �   |   ~   �      d            " Computed Q=" & to_hstring(unsigned(ho)) & ", Expected Q=" & to_hstring(unsigned(Hov)) 5��    |   c                                       5�_�   �   �           �   v       ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f٦     �   u   w   �      h            " Computed Q=" & to_hstring(unsigned(ao)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    u                     �                     5�_�   �   �           �   w       ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f٨     �   v   x   �      h            " Computed Q=" & to_hstring(unsigned(bo)) & ", Expected Q=" & to_hstring(unsigned(Bov)) &LF&5��    v                     @                     5�_�   �   �           �   x       ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f٩     �   w   y   �      h            " Computed Q=" & to_hstring(unsigned(co)) & ", Expected Q=" & to_hstring(unsigned(Cov)) &LF&5��    w                     �                     5�_�   �   �           �   y       ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f٪     �   x   z   �      h            " Computed Q=" & to_hstring(unsigned(do)) & ", Expected Q=" & to_hstring(unsigned(Dov)) &LF&5��    x                                          5�_�   �   �           �   z       ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f٫     �   y   {   �      h            " Computed Q=" & to_hstring(unsigned(eo)) & ", Expected Q=" & to_hstring(unsigned(Eov)) &LF&5��    y                     ~                     5�_�   �   �           �   {       ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    f٭     �   z   |   �      h            " Computed Q=" & to_hstring(unsigned(fo)) & ", Expected Q=" & to_hstring(unsigned(Fov)) &LF&5��    z                     �                     5�_�   �   �           �   |       ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    fٯ     �   {   }   �      h            " Computed Q=" & to_hstring(unsigned(go)) & ", Expected Q=" & to_hstring(unsigned(Gov)) &LF&5��    {                     R                     5�_�   �               �   }       ����                                                                                                                                                                                                                                                                                                                            ~          ~   5       v   5    fٰ   
 �   |   ~   �      c            " Computed Q=" & to_hstring(unsigned(ho)) & ", Expected Q=" & to_hstring(unsigned(Hov))5��    |                     �                     5�_�   �           �   �   v       ����                                                                                                                                                                                                                                                                                                                            x          x   5       v   5    f�D     �   v   w   �    �   v   w   �      h            " Computed Q=" & to_hstring(unsigned(ao)) & ", Expected Q=" & to_hstring(unsigned(Aov)) &LF&5��    v                      2              i       5�_�   �   �       �   �   v   6    ����                                                                                                                                                                                                                                                                                                                            s          u          V       e��1     �   u   w   �      A            " Computed Q=" & integer'image(to_integer((ao))) &LF&5��    u   6                  �                     5�_�   �   �           �   v   6    ����                                                                                                                                                                                                                                                                                                                            s          u          V       e��3     �   u   w   �      @            " Computed Q=" & integer'image(to_integer(ao))) &LF&5��    u   6                  �                     5�_�   �   �           �   v   8    ����                                                                                                                                                                                                                                                                                                                            s          u          V       e��4     �   u   w   �      ?            " Computed Q=" & integer'image(to_integer(ao)) &LF&5��    u   8                  �                     5�_�   �   �           �   w   6    ����                                                                                                                                                                                                                                                                                                                            s          u          V       e��5     �   v   x   �      =            " Expected Q=" & integer'image(to_integer((Aov)))5��    v   6                  ;                     5�_�   �   �           �   w   6    ����                                                                                                                                                                                                                                                                                                                            s          u          V       e��6     �   v   x   �      <            " Expected Q=" & integer'image(to_integer(Aov)))5��    v   6                  ;                     5�_�   �   �           �   w   9    ����                                                                                                                                                                                                                                                                                                                            s          u          V       e��6     �   v   x   �      ;            " Expected Q=" & integer'image(to_integer(Aov))5��    v   9                  >                     5�_�   �   �   �       �   w   :    ����                                                                                                                                                                                                                                                                                                                            s          u          V       e��P     �   v   x   �      :            " Expected Q=" & integer'image(to_integer(Aov)5��    v   :                  ?                     5�_�   �               �   w   :    ����                                                                                                                                                                                                                                                                                                                            s          u          V       e��V    �   v   x   �      ;            " Expected Q=" & integer'image(to_integer(Aov))5��    v   :                  ?                     5�_�   �           �   �   w   6    ����                                                                                                                                                                                                                                                                                                                            s          u          V       e��J     �   v   x        5��    v                            <               5�_�   �       �   �   �      	    ����                                                                                                                                                                                                                                                                                                                            r          t          V       e���     �              5��                                                5�_�   �           �   �      	    ����                                                                                                                                                                                                                                                                                                                            r          t          V       e���     �              5��                          "                      5�_�   �           �   �   s       ����                                                                                                                                                                                                                                                                                                                            V          W          V       e��     �   r   t   �      <            " =" & integer'image(to_integer(signed(x))) &LF&5��    r                                          5�_�   z           |   {   \        ����                                                                                                                                                                                                                                                                                                                            V          W          V       e�ߋ     �   \   ]   p    �   \   ]   p                  read(tb_line, Aov);   !            read(tb_line, space);5��    \                      �
              B       5�_�   I           K   J   0       ����                                                                                                                                                                                                                                                                                                                                                       e�ޕ     �   0   1   g    �   0   1   g      :        variable Xv, Yv, Zv, res: bit_vector(31 downto 0);5��    0                      h              ;       5�_�   .   0       3   /   !       ����                                                                                                                                                                                                                                                                                                                                                V       e��     �   !   "   `    �   !   "   `                        hi => hi, 5��    !                      S                     5�_�   /   1           0   "       ����                                                                                                                                                                                                                                                                                                                                                V       e��     �   "   #   a    �   "   #   a                        hi => hi, 5��    "                      p                     5�_�   0   2           1   #       ����                                                                                                                                                                                                                                                                                                                                                V       e��     �   #   $   b    �   #   $   b                        hi => hi, 5��    #                      �                     5�_�   1               2   $       ����                                                                                                                                                                                                                                                                                                                                                V       e��     �   $   %   c    �   $   %   c                        hi => hi, 5��    $                      �                     5�_�                            ����                                                                                                                                                                                                                                                                                                                            4          6          V       e��0     �         ^                        i => ci, 5��                         �                     5�_�             
             ����                                                                                                                                                                                                                                                                                                                            ,          .          V       e��K     �          V      :        variable Av, Yv, Zv, res: bit_vector(31 downto 0);5��                        �                    5�_�      	                     ����                                                                                                                                                                                                                                                                                                                            ,          .          V       e��R     �          V      :        variable Av, Bv, Zv, res: bit_vector(31 downto 0);5��                        �                    5�_�                  	          ����                                                                                                                                                                                                                                                                                                                            ,          .          V       e��V     �          V      :        variable Av, Bv, uv, res: bit_vector(31 downto 0);5��                        �                    5��