Vim�UnDo� �/u|���M<�P���[����Y��.:D��   �                Q      Q  Q  Q    f)#�    _�                             ����                                                                                                                                                                                                                                                                                                                                                             f'�z     �                   �               5��                                          �       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'�|     �                 end sha256_1b ;5��                         �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'ׁ     �                e n t i t y sha256_1b i s5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'ׁ     �                en t i t y sha256_1b i s5��                                                5�_�                          ����                                                                                                                                                                                                                                                                                                                                                             f'ׄ     �                ent i t y sha256_1b i s5��                                                5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                             f'ׅ     �                enti t y sha256_1b i s5��                                                5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                             f'ׅ     �                entit y sha256_1b i s5��                                                5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                             f'׈     �                entity sha256_1b i s5��                                                5�_�   
                         ����                                                                                                                                                                                                                                                                                                                                                             f'׉     �               po r t (5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'׋     �                   po r t (5��                                               5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'׋     �                   por t (5��                                               5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f'׍     �               clock , r e s e t : in b i t ;5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'׏     �               &        clock , r e s e t : in b i t ;5��                         0                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'׏     �               %        clock , re s e t : in b i t ;5��                         1                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'׏     �               $        clock , res e t : in b i t ;5��                         2                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'א     �               #        clock , rese t : in b i t ;5��                         3                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'ג     �               "        clock , reset : in b i t ;5��                         ;                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'ג     �               !        clock , reset : in bi t ;5��                         <                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'ד     �                        clock , reset : in bit ;5��                         =                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f'ה     �               s e r i a l _ i n : in b i t ;5��                          ?                      5�_�                       	    ����                                                                                                                                                                                                                                                                                                                                                             f'ו     �               &        s e r i a l _ i n : in b i t ;5��       	                  H                      5�_�                       
    ����                                                                                                                                                                                                                                                                                                                                                             f'ז     �               %        se r i a l _ i n : in b i t ;5��       
                  I                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'ז     �               $        ser i a l _ i n : in b i t ;5��                         J                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'ז     �               #        seri a l _ i n : in b i t ;5��                         K                      5�_�      !                     ����                                                                                                                                                                                                                                                                                                                                                             f'ז     �               "        seria l _ i n : in b i t ;5��                         L                      5�_�      "          !          ����                                                                                                                                                                                                                                                                                                                                                             f'ך     �               !        serial _ i n : in b i t ;5��                         M                      5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                                                             f'ך     �                        serial_ i n : in b i t ;5��                         N                      5�_�   "   $           #          ����                                                                                                                                                                                                                                                                                                                                                             f'כ     �                       serial_i n : in b i t ;5��                         O                      5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                                             f'ל     �                       serial_in : in b i t ;5��                         W                      5�_�   $   &           %          ����                                                                                                                                                                                                                                                                                                                                                             f'ם     �                       serial_in : in bi t ;5��                         X                      5�_�   %   '           &          ����                                                                                                                                                                                                                                                                                                                                                             f'ם     �                       serial_in : in bit ;5��                         Y                      5�_�   &   (           '           ����                                                                                                                                                                                                                                                                                                                                                             f'מ     �               s e r i a l _ o u t : out b i t5��                          [                      5�_�   '   )           (      	    ����                                                                                                                                                                                                                                                                                                                                                             f'נ     �               '        s e r i a l _ o u t : out b i t5��       	                  d                      5�_�   (   *           )      
    ����                                                                                                                                                                                                                                                                                                                                                             f'נ     �               &        se r i a l _ o u t : out b i t5��       
                  e                      5�_�   )   +           *          ����                                                                                                                                                                                                                                                                                                                                                             f'נ     �               %        ser i a l _ o u t : out b i t5��                         f                      5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                                             f'ס     �               $        seri a l _ o u t : out b i t5��                         g                      5�_�   +   -           ,          ����                                                                                                                                                                                                                                                                                                                                                             f'ס     �               #        seria l _ o u t : out b i t5��                         h                      5�_�   ,   .           -          ����                                                                                                                                                                                                                                                                                                                                                             f'ס     �               "        serial _ o u t : out b i t5��                         i                      5�_�   -   /           .          ����                                                                                                                                                                                                                                                                                                                                                             f'ס     �               !        serial_ o u t : out b i t5��                         j                      5�_�   .   0           /          ����                                                                                                                                                                                                                                                                                                                                                             f'ע     �                        serial_o u t : out b i t5��                         k                      5�_�   /   1           0          ����                                                                                                                                                                                                                                                                                                                                                             f'ע     �                       serial_ou t : out b i t5��                         l                      5�_�   0   2           1          ����                                                                                                                                                                                                                                                                                                                                                             f'פ     �                       serial_out : out b i t5��                         u                      5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                                                             f'פ     �                       serial_out : out bi t5��                         v                      5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                                                             f'צ     �                       serial_out : out bit5��                         m                      5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                                                             f'ק     �                       serial_in : in bit;5��                         P                      5�_�   4   6           5           ����                                                                                                                                                                                                                                                                                                                                                             f'ש    �               ) ;5��                          v                      5�_�   5   7           6           ����                                                                                                                                                                                                                                                                                                                                                             f(J�     �                 end architecture �      
         architecture rtl of  is�                     �                 arch�                  �               5��                          �                      �                          �                      �                          �                      �                         �                      �                         �                     �                         �                     �                         �                     �                         �                     �                        �                      �                          �                       �                        �                      �                         �                      �                         �                      �                         �                      5�_�   6   8           7   	       ����                                                                                                                                                                                                                                                                                                                            	          	          v       f(J�     �   	   
       �                 end architecture rtl;�   	   
       �   	   
       �   	   
       �   	   
       �   	   
       �   	   
       �   	   
       �   	   
       �   	   
       �      
         architecture rtl of sha256 is5��                        �                     �                        �                     �                         �                      �                        �                     �                         �                      �                        �                     �                         �                      �                        �                     �                         �                      �                        �                     �                         �                      �                        �                     �                         �                      �                        �                     �                         �                      �                        �                     �                         �                      �                     	   �              	       �                         �                      �              	       
   �       	       
       5�_�   7   9           8   	       ����                                                                                                                                                                                                                                                                                                                            	           	          v       f(J�    �      
         $architecture Behavioral of sha256 is5��                        �                     �                        �                     �                         �                      �                         �                      �                     	   �              	       �              	          �       	              �                     	   �              	       5�_�   8   :           9           ����                                                                                                                                                                                                                                                                                                                                                             f(m�     �      S       �             5��                   E       �               �	      5�_�   9   ;           :          ����                                                                                                                                                                                                                                                                                                                                                             f(m�     �                    5��                          �                      5�_�   :   <           ;   	       ����                                                                                                                                                                                                                                                                                                                                                             f(ӹ     �   	      T          �   	      S    5��    	                      �                      �    	                      �                      �    	                      �                      �    	                     �                      �    
                     �                      5�_�   ;   =           <          ����                                                                                                                                                                                                                                                                                                                                                             f(��     �         U    �         U    5��                          �                      5�_�   <   ?           =          ����                                                                                                                                                                                                                                                                                                                                                             f(��     �         V          signal sender_clk: bit;5��                        �                     5�_�   =   @   >       ?          ����                                                                                                                                                                                                                                                                                                                                                             f(��     �         V    �         V    5��                          �                      5�_�   ?   A           @          ����                                                                                                                                                                                                                                                                                                                                                             f(��     �         W          signal receiver_clk: bit;5��                        �                     5�_�   @   B           A   
        ����                                                                                                                                                                                                                                                                                                                                                             f(�0     �   	      W    5��    	                      �                      �    	                      �                      �    	                      �                      5�_�   A   C           B   
        ����                                                                                                                                                                                                                                                                                                                                                             f(�1     �   
      X    �   
      X    5��    
               	       �               �       5�_�   B   D           C          ����                                                                                                                                                                                                                                                                                                                                                             f(�?     �         d              generic�         c          send_clk: sender_clk�         b          �         a    5��                          �                     �                          �                     �                          �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                     
   �             
       �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                     
   �             
       �              
          �      
              �                     
   �             
       �                        �                     �                         �                     �                        �                    �                        �                    �                        �                    5�_�   C   E           D          ����                                                                                                                                                                                                                                                                                                                                                             f(�[     �         d              generic map5��                         �                     5�_�   D   F           E          ����                                                                                                                                                                                                                                                                                                                                                             f(�]     �         e              port�         d              generic map()5��                        �              	       �                         �                     �                        �                    �                        �                    �                        �                    5�_�   E   G           F          ����                                                                                                                                                                                                                                                                                                                                                             f(�_     �         e              port map5��                         �                     5�_�   F   H           G          ����                                                                                                                                                                                                                                                                                                                                                             f(�b     �         e              port map()5��                         �                     5�_�   G   I           H          ����                                                                                                                                                                                                                                                                                                                                                             f(�e     �         e              port map(clock)5��                                              �                     
                
       �              
                
              �                     
                
       5�_�   H   J           I      #    ����                                                                                                                                                                                                                                                                                                                                                             f(�i     �         e      #        port map(clock, sender_clk)5��       #                                       5�_�   I   K           J           ����                                                                                                                                                                                                                                                                                                                                         #       V   #    f(�m     �         e    5��                                        	       �                                               5�_�   J   L           K           ����                                                                                                                                                                                                                                                                                                                                         #       V   #    f(�n     �      "   f    �         f    5��                                        T       5�_�   K   M           L   !       ����                                                                                                                                                                                                                                                                                                                                         #       V   #    f(�o     �   !   #   i    5��    !                      g              	       �    !                      g                     5�_�   L   O           M   "        ����                                                                                                                                                                                                                                                                                                                                         #       V   #    f(�p     �   "   &   j    �   "   #   j    5��    "                      h              T       5�_�   M   P   N       O           ����                                                                                                                                                                                                                                                                                                                                      !          V       f(Ԑ     �       "          $        port map(clock, sender_clk);�          m          send_clk: sender_clk5��                                            �                        $                    �                         `                    5�_�   O   Q           P          ����                                                                                                                                                                                                                                                                                                                                      !          V       f(ԕ     �          m          receive_clk: receiveer_clk5��                         *                     5�_�   P   R           Q   !       ����                                                                                                                                                                                                                                                                                                                                      !          V       f(Ԙ     �       "   m      '        port map(clock, receiveer_clk);5��                          f                     5�_�   Q   S           R          ����                                                                                                                                                                                                                                                                                                                                      !          V       f(ԥ     �          m          receive_clk: receiver_clk5��                        $                    5�_�   R   T           S          ����                                                                                                                                                                                                                                                                                                                                      !          V       f(Ԫ     �         m          send_clk: sender_clk5��              
          �      
              �                         �                     �                         �                     �                         �                     �                        �                    �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    5�_�   S   U           T   #        ����                                                                                                                                                                                                                                                                                                                                      !          V       f(Լ     �   "   #              send_clk: sender_clk           generic map()   $        port map(clock, sender_clk);       5��    "                      i      Y               5�_�   T   V           U          ����                                                                                                                                                                                                                                                                                                                                      !          V       f(��     �         j          �         i    5��                          �                     �                         �                     5�_�   U   W           V          ����                                                                                                                                                                                                                                                                                                                                       "          V       f(�     �         j              generic map()5��                                               5�_�   V   X           W          ����                                                                                                                                                                                                                                                                                                                                       "          V       f(�     �         j              generic map(2)5��                                              �       +                                       5�_�   W   Y           X   "   %    ����                                                                                                                                                                                                                                                                                                                                       "   &       V   *    f(��     �      #   j          receive_clk: slow_clk           generic map()   &        port map(clock, receiver_clk);5��                         >      W       `       5�_�   X   Z           Y   "   %    ����                                                                                                                                                                                                                                                                                                                                       "   &       V   *    f(��     �   "   $   k              �   "   $   j    5��    "                      �                     �    "                     �                    �    "                    �                    �    "                     �                     �    "                     �                     �    "                     �                     �    "                    �                    �    "                    �                    �    "                    �                    �    "                     �                     �    "                     �                     �    "                    �                    �    "                    �                    �    "                    �                    5�_�   Y   [           Z   #       ����                                                                                                                                                                                                                                                                                                                                       "   &       V   *    f(��     �   "   $   k          receiver_clk <= clock5��    "                     �                     5�_�   Z   \           [          ����                                                                                                                                                                                                                                                                                                                                       "   &       V   *    f(��     �                    signal encrypt_clk: bit;5��                          �                     5�_�   [   ]           \   "       ����                                                                                                                                                                                                                                                                                                                                      !   &       V   *    f(��     �   !   "              receiver_clk <= clock;5��    !                      �                     5�_�   \   ^           ]           ����                                                                                                                                                                                                                                                                                                                                      !   &       V   *    f(��     �          i    �          i    5��                          !                     5�_�   ]   _           ^          ����                                                                                                                                                                                                                                                                                                                                       "   &       V   *    f(��     �         j          send_clk: slow_clk5��                      
   �              
       5�_�   ^   `           _          ����                                                                                                                                                                                                                                                                                                                                       "   &       V   *    f(�      �         j              clock , reset : in bit;5��                         >                      5�_�   _   a           `           ����                                                                                                                                                                                                                                                                                                                                       "   &       V   *    f(�     �         j           send_clk: slow_clk -- Envia 5��                          �                     �                         �                    5�_�   `   b           a          ����                                                                                                                                                                                                                                                                                                                                       "   &       V   *    f(�     �          j          receiver_clk <= clock;5��                         ^                     5�_�   a   c           b      )    ����                                                                                                                                                                                                                                                                                                                                       "   &       V   *    f(�#     �          j      )    receiver_clk <= clock; -- recebe a 5k5��       )                  m                     5�_�   b   d           c   $       ����                                                                                                                                                                                                                                                                                                                                       "   &       V   *    f(�B     �   #   %   j          process(new_clk) is5��    #                    �                    5�_�   c   e           d   $       ����                                                                                                                                                                                                                                                                                                                                       "   &       V   *    f(�T     �   #   %   j          process(clock) is5��    #                     �                     5�_�   d   f           e   &       ����                                                                                                                                                                                                                                                                                                                                       "   &       V   *    f(�Y     �   %   '   j      $        if rising_edge(new_clk) then5��    %                    '                    5�_�   e   g           f          ����                                                                                                                                                                                                                                                                                                                                       "   &       V   *    f(�v     �         j    5��                          �                     �                          �                     5�_�   f   h           g           ����                                                                                                                                                                                                                                                                                                                            !          #   &       V   *    f(�v     �         k    �         k    5��                          �              �       5�_�   g   i           h      	    ����                                                                                                                                                                                                                                                                                                                            #          %   &       V   *    f(�x     �         m      ;    type transmiter is (starting, sending, stopping, idle);5��       	       
          �      
              �                         �                     �       
                  �                     �       	              	   �             	       5�_�   h   j           i          ����                                                                                                                                                                                                                                                                                                                            #          %   &       V   *    f(ׇ     �         m      L    signal state: transmiter := idle; -- Declaração da máquina de estados5��              
          �      
              �                         �                     �                         �                     �                     	   �             	       �              	       	   �      	       	       �              	          �      	              �                     	   �             	       5�_�   i   k           j          ����                                                                                                                                                                                                                                                                                                                            #          %   &       V   *    f(א     �         m      :    type sha_state is (starting, sending, stopping, idle);5��                        �                    �                        �                    5�_�   j   l           k      +    ����                                                                                                                                                                                                                                                                                                                            #          %   &       V   *    f(ט     �         m      ;    type sha_state is (receiving, sending, stopping, idle);5��       +                 �                    5�_�   k   m           l      +    ����                                                                                                                                                                                                                                                                                                                            #          %   &       V   *    f(ל     �         m      ;    type sha_state is (receiving, sending, mutating, idle);5��       +                 �                    5�_�   l   n           m          ����                                                                                                                                                                                                                                                                                                                            #          %   &       V   *    f(ض     �   
      m    5��    
                      �                      �    
                      �                      5�_�   m   o           n           ����                                                                                                                                                                                                                                                                                                                            $          &   &       V   *    f(ط     �   
      o          �   
      n    5��    
                      �                      �    
                   
   �               
       �    
   	                  �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                 	   �              	       �    
          	          �       	              �    
                    �                     �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                 
   �              
       �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                 	   �              	       �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                 	   �              	       �    
          	          �       	              �    
                 	   �              	       5�_�   n   p           o          ����                                                                                                                                                                                                                                                                                                                            %          '   &       V   *    f(ؾ     �         p          end component�   
      o          component serial_in5��    
                    �                      �                         �                     �                         �                     �                         �                      �                         �                      �       
                  �                      �       	                  �                      �                     	   �              	       �              	          �       	              �                     
   �              
       5�_�   o   q           p          ����                                                                                                                                                                                                                                                                                                                            &          (   &       V   *    f(��     �         p    �         p    5��                          �               �       5�_�   p   r           q          ����                                                                                                                                                                                                                                                                                                                                                       f(��     �         x              WIDTH: natural := 7       );   	    port(   *        clock, reset, serial_data: in bit;   "        done, parity_bit: out bit;   7        parallel_data: out bit_vector(WIDTH-1 downto 0)       );�         x          generic(5��                         �                      �                         �                      �                                              �                         $                     �                         2                     �                         a                     �                         �                     �                         �                     5�_�   q   s           r          ����                                                                                                                                                                                                                                                                                                                                                       f(��     �   
      x          component serial_in5��    
          	          �       	              5�_�   r   t           s   7       ����                                                                                                                                                                                                                                                                                                                                                       f(�	     �   6   8   x                      done <= '1';5��    6                    '                    �    6                     )                     �    6                     (                     �    6                 	   '             	       �    6                     /                     �    6                     .                     �    6                     -                     �    6                     ,                     �    6                     +                     �    6                     *                     �    6                     )                     �    6                     (                     �    6                    '                    �    6                     1                     �    6                     0                     �    6                     /                     �    6                     .                     �    6                     -                     �    6                     ,                     �    6                     +                     �    6                     *                     �    6                     )                     �    6                     (                     �    6                 
   '             
       �    6          
       
   '      
       
       �    6          
          '      
              �    6                 
   '             
       5�_�   s   u           t   9        ����                                                                                                                                                                                                                                                                                                                            9          <          V       f(�     �   8   9                          -- Control   $                start_signal <= '0';   "                start_stop <= '0';   "                shift_data <= '0';5��    8                      ;      �               5�_�   t   v           u   =       ����                                                                                                                                                                                                                                                                                                                            =          =   ;       v   ;    f(�&     �   <   >   t      A                        if start = '1' and serial_data = '0' then5��    <          !          �      !              �    <                     �                     �    <                     �                     �    <                 
   �             
       �    <          
       	   �      
       	       �    <   #                  �                     5�_�   u   w           v   =       ����                                                                                                                                                                                                                                                                                                                            =          =   ;       v   ;    f(�B     �   <   >   t      (                        if serial_i then5��    <                    �                    �    <                     �                     �    <                     �                     �    <                 
   �             
       �    <          
          �      
              �    <                 
   �             
       �    <   $                  �                     �    <   #                  �                     �    <   "                 �                    5�_�   v   x           w   =   '    ����                                                                                                                                                                                                                                                                                                                            =          =   ;       v   ;    f(�G     �   <   >   t      ,                        if serial_in =  then5��    <   '                  �                     5�_�   w   y           x   =   (    ����                                                                                                                                                                                                                                                                                                                            =          =   ;       v   ;    f(�G     �   <   >   t      .                        if serial_in = '' then5��    <   (                  �                     5�_�   x   z           y   >   %    ����                                                                                                                                                                                                                                                                                                                            =          =   ;       v   ;    f(�J     �   =   ?   t      .                            state <= starting;5��    =   %                 �                    �    =   (                  �                     �    =   '                  �                     �    =   &                  �                     �    =   %                 �                    �    =   0                  �                     �    =   /                  �                     �    =   .                  �                     �    =   -                  �                     �    =   ,                  �                     �    =   +                  �                     �    =   *                  �                     �    =   )                  �                     �    =   (                  �                     �    =   '                  �                     �    =   &                  �                     �    =   %                 �                    �    =   *                  �                     �    =   )                  �                     �    =   (                  �                     �    =   '                  �                     �    =   &                  �                     �    =   %                 �                    �    =   ,                  �                     �    =   +                  �                     �    =   *                  �                     �    =   )                  �                     �    =   (                  �                     �    =   '                  �                     �    =   &                  �                     �    =   %              	   �             	       �    =   %       	       	   �      	       	       �    =   %       	          �      	              �    =   %              	   �             	       5�_�   y   {           z   ?   '    ����                                                                                                                                                                                                                                                                                                                            =          =   ;       v   ;    f(�U     �   >   ?          (                            done <= '0';5��    >                      �      )               5�_�   z   |           {   A        ����                                                                                                                                                                                                                                                                                                                            =          =   ;       v   ;    f(�W     �   @   A          0                            start_signal <= '1';5��    @                            1               5�_�   {   }           |   A        ����                                                                                                                                                                                                                                                                                                                            =          =   ;       v   ;    f(�W     �   @   A          .                            shift_data <= '1';5��    @                            /               5�_�   |   ~           }   @        ����                                                                                                                                                                                                                                                                                                                            =          =   ;       v   ;    f(�X     �   ?   @          &                            -- Control5��    ?                      �      '               5�_�   }              ~   0        ����                                                                                                                                                                                                                                                                                                                            =          =   ;       v   ;    f(�_     �   2   4   s              generic�   1   4   r          receiver�   0   3   q          �   0   2   p    5��    0                      �                     �    0                      �                     �    0                     �                     �    1                     �                     �    1                     �                     �    1                     �                     �    1                     �                     �    1                     �                     �    1                    �                    �    1                    �                    �    1                    �                    �    1                     �                     �    1                     �                     �    1                    �                    �    1                    �                    �    1                     �                     �    1                     �                     �    1                     �                     �    1                    �                    �    1                    �                    �    1                    �                    �    1                     �                     �    2                     �                     �    2                    �                    �    2                    �                    �    2                    �                    5�_�   ~   �              3       ����                                                                                                                                                                                                                                                                                                                            @          @   ;       v   ;    f(�|     �   2   4   s              generic map5��    2                     �                     5�_�      �           �   3       ����                                                                                                                                                                                                                                                                                                                            @          @   ;       v   ;    f(�~     �   2   4   s              generic map()5��    2                     �                     5�_�   �   �           �   3       ����                                                                                                                                                                                                                                                                                                                            @          @   ;       v   ;    f(ـ     �   3   5   t              port�   2   5   s              generic map(8)5��    2                    �              	       �    3                     �                     �    3                    �                    �    3                    �                    �    3                    �                    5�_�   �   �           �   4       ����                                                                                                                                                                                                                                                                                                                            A          A   ;       v   ;    f(ق     �   3   5   t              port map5��    3                     �                     5�_�   �   �           �   4       ����                                                                                                                                                                                                                                                                                                                            A          A   ;       v   ;    f(ل     �   3   6   u              port map(�   4   6                          )�   3   6   t              port map()5��    3                    �              	       �    4                     �                    �    3                    �              	       �    4                     �                     �    4                      �                     5�_�   �   �           �   6       ����                                                                                                                                                                                                                                                                                                                            C          C   ;       v   ;    f(ه     �   5   7   v                      )5��    5                     �                     5�_�   �   �           �   6   	    ����                                                                                                                                                                                                                                                                                                                            C          C   ;       v   ;    f(ى     �   5   7   v      	        )5��    5   	                  �                     5�_�   �   �           �   5        ����                                                                                                                                                                                                                                                                                                                            C          C   ;       v   ;    f(ي     �   4   6   v       5��    4                      �                     �    4                    �                    �    4                    �                    �    4                    �                    �    4                    �                    �    4                     �                     �    4                     �                     �    4                     �                     �    4                 	   �             	       �    4                     �                     �    4                     �                     �    4                     �                     �    4                     �                     �    4                     �                     �    4                     �                     �    4                     �                     �    4                     �                     �    4                    �                    �    4                    �                    �    4                    �                    �    4                    �                    5�_�   �   �           �   5   !    ����                                                                                                                                                                                                                                                                                                                            C          C   ;       v   ;    f(ٛ     �   6   8   x                  serial_data�   5   8   w                  reset�   4   7   v      !            clock => receiver_clk5��    4   !                  �                     �    4   "                 �                     �    5                     �                     �    5                    �                    �    5                    �                    �    5                    �                    �    5                                        �    5                                         �    6                                          �    6                                        �    6                                        �    6                                        �    6                                        �    6                 
                
       �    6          
       	         
       	       �    6          	       	         	       	       �    6          	                	              �    6                 	                	       5�_�   �   �           �   7   $    ����                                                                                                                                                                                                                                                                                                                            E          E   ;       v   ;    f(ٸ     �   6   9   x      $            serial_data => serial_in5��    6   $                  '                     �    6   %                 (                     �    7                     5                     5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            F          F   ;       v   ;    f(��     �   $   &   y    5��    $                      D                     5�_�   �   �           �   %        ����                                                                                                                                                                                                                                                                                                                            G          G   ;       v   ;    f(��     �   $   (   z          5��    $                     D                    �    %                      E                     �    %                    Y                    �    %                    [                     �    &                     `                     5�_�   �   �           �   ;       ����                                                                                                                                                                                                                                                                                                                            I          I   ;       v   ;    f(��     �   :   =   |                  done =>5��    :                     x                     �    :                    y                    �    :                    y                    �    :                    y                    �    :   '                 �                     �    ;                      �                     5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            J          J   ;       v   ;    f(�
     �   $   (   ~          �   $   &   }    5��    $                      D                     �    $                      D                     �    $                     D                     �    %                     I                     �    %                    P                     �    &                     U                     �    &                     a                     �    &                     `                     �    &                     _                     �    &                     ^                     �    &                     ]                     �    &                     \                     �    &   
                 [                    5�_�   �   �           �   ?        ����                                                                                                                                                                                                                                                                                                                            M          M   ;       v   ;    f(�      �   >   @   �       5��    >                      �                     �    >                    �                    �    >                    �                    �    >                    �                    �    >          	          �      	              �    >                    �                    �    >                    �                    �    >                    �                    5�_�   �   �           �   ?       ����                                                                                                                                                                                                                                                                                                                            M          M   ;       v   ;    f(�+     �   >   A   �                  data_parity5��    >                     �                     �    >                    �                     �    ?                      �                     5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            N          N   ;       v   ;    f(�9     �   '   )   �          �   '   )   �    5��    '                      n                     �    '                     r                     �    '                     �                     �    '                     �                     �    '                     �                     �    '                     �                     �    '                 
   �             
       �    '          
          �      
              �    '                 
   �             
       5�_�   �   �           �   (   $    ����                                                                                                                                                                                                                                                                                                                            O          O   ;       v   ;    f(�[     �   '   )   �      $    signal received_data: bit_vector5��    '   $                  �                     5�_�   �   �           �   (   %    ����                                                                                                                                                                                                                                                                                                                            O          O   ;       v   ;    f(�\     �   '   )   �      &    signal received_data: bit_vector()5��    '   %                  �                     �    '   '                 �                    �    '   '                 �                    �    '   '              	   �             	       �    '   /                  �                     5�_�   �   �           �   (   0    ����                                                                                                                                                                                                                                                                                                                            O          O   ;       v   ;    f(�`     �   '   )   �      0    signal received_data: bit_vector(7 downto 0)5��    '   0                  �                     5�_�   �   �           �   A        ����                                                                                                                                                                                                                                                                                                                            O          O   ;       v   ;    f(�d     �   @   B   �       5��    @                                           �    @                 
                
       �    @          
                
              �    @                                        �    @                                        �    @                                        �    @                                        �    @                                        �    @                                        5�_�   �   �           �   J        ����                                                                                                                                                                                                                                                                                                                            O          O   ;       v   ;    f(��     �   J   L   �                      �   J   L   �    5��    J                      �                     �    J                      �                     �    J                                        �    J                                        �    J                                        5�_�   �   �           �   K   &    ����                                                                                                                                                                                                                                                                                                                            P          P   ;       v   ;    f(��     �   J   L   �      &                finished_receiving <= 5��    J   &                                       5�_�   �   �           �   K   '    ����                                                                                                                                                                                                                                                                                                                            P          P   ;       v   ;    f(��     �   J   L   �      (                finished_receiving <= ''5��    J   '                                       5�_�   �   �           �   K   )    ����                                                                                                                                                                                                                                                                                                                            P          P   ;       v   ;    f(��     �   J   L   �      )                finished_receiving <= '0'5��    J   )                                       5�_�   �   �           �   K   '    ����                                                                                                                                                                                                                                                                                                                            P          P   ;       v   ;    f(��     �   J   L   �      *                finished_receiving <= '0';5��    J   '                                     5�_�   �   �           �   K   '    ����                                                                                                                                                                                                                                                                                                                            P          P   ;       v   ;    f(��     �   J   K          *                finished_receiving <= '1';5��    J                      �      +               5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            O          O   ;       v   ;    f(�     �   S   U   �      $                    when starting =>5��    S                    �                    �    S                    �                    �    S                 	   �             	       �    S          	       	   �      	       	       �    S          	          �      	              �    S                 	   �             	       5�_�   �   �           �   T        ����                                                                                                                                                                                                                                                                                                                            O   !       R          V   !    f(�
     �   T   Y   �    �   T   U   �    5��    T                      �              �       5�_�   �   �   �       �   U       ����                                                                                                                                                                                                                                                                                                                            O   !       R          V   !    f(�     �   T   V   �      /                        if serial_in = '0' then5��    T          	                	              �    T                                        �    T                                        �    T                                        5�_�   �   �           �   U   1    ����                                                                                                                                                                                                                                                                                                                            O   !       R          V   !    f(�;     �   T   V   �      8                        if finished_receiving = '0' then5��    T   1                                     5�_�   �   �           �   V   %    ����                                                                                                                                                                                                                                                                                                                            O   !       R          V   !    f(�A     �   U   W   �      /                            state <= receiving;5��    U   %       	          H      	              �    U   %                 H                    �    U   %                 H                    �    U   %                 H                    5�_�   �   �           �   V   ,    ����                                                                                                                                                                                                                                                                                                                            O   !       R          V   !    f(�G     �   U   W   �      -                            state <= encrypt;5��    U   ,                  O                     5�_�   �   �           �   #   2    ����                                                                                                                                                                                                                                                                                                                            O   !       R          V   !    f(�N     �   "   $   �      :    type sha_state is (receiving, sending, encrypt, idle);5��    "   2                  �                     5�_�   �   �           �   Y   (    ����                                                                                                                                                                                                                                                                                                                            O   !       R          V   !    f(�Y     �   X   Y          )                        state <= sending;   ,                        start_signal <= '0';5��    X                      x      W               5�_�   �   �           �   M        ����                                                                                                                                                                                                                                                                                                                            O   !       R          V   !    f(�]     �   L   M           5��    L                      #                     5�_�   �   �   �       �   X        ����                                                                                                                                                                                                                                                                                                                            S           W           V        f(�l     �   X   ^   �    �   X   Y   �    5��    X                      x              �       5�_�   �   �           �   ]       ����                                                                                                                                                                                                                                                                                                                            S           W           V        f(�n     �   ]   _   �    5��    ]                      )	                     �    ]                      )	                     5�_�   �   �           �   Y       ����                                                                                                                                                                                                                                                                                                                            S           W           V        f(�r     �   X   Z   �      %                    when receiving =>5��    X          	          �      	              �    X                 
   �             
       �    X          
          �      
              �    X                 
   �             
       5�_�   �   �           �   B   	    ����                                                                                                                                                                                                                                                                                                                            S           W           V        f(��     �   B   F   �              �   B   D   �    5��    B                      ;              	       �    B                      ;                     �    B                     ;              	       �    C                    @                    �    C                    @                    �    C                    S                     �    D                     X                     5�_�   �   �           �   E       ����                                                                                                                                                                                                                                                                                                                            V           Z           V        f(��     �   D   F   �              port map5��    D                     d                     5�_�   �   �           �   E       ����                                                                                                                                                                                                                                                                                                                            V           Z           V        f(�     �   D   G   �              port map(�   E   G                          )�   D   G   �              port map()5��    D                    e              	       �    E                     f                    �    D                    e              	       �    E                      f                     5�_�   �   �           �   G       ����                                                                                                                                                                                                                                                                                                                            X           \           V        f(�     �   F   H   �                      )5��    F                     o                     5�_�   �   �           �   G   	    ����                                                                                                                                                                                                                                                                                                                            X           \           V        f(�     �   F   H   �      	        )5��    F   	                  p                     5�_�   �   �           �   F        ����                                                                                                                                                                                                                                                                                                                            X           \           V        f(�	     �   E   I   �       5��    E                      f                     �    E                    x                     �    F                     �                     �    F                    �                     �    G                     �                     5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                            Z           ^           V        f(�"     �   (   *   �          �   (   *   �    5��    (                      �                     �    (                     �                     �    (                    �                    �    (                 
   �             
       �    (          
       
   �      
       
       �    (          
          �      
              �    (                    �                    �    (   !                  �                     5�_�   �   �           �   )   !    ����                                                                                                                                                                                                                                                                                                                            [           _           V        f(�.     �   (   *   �      !    signal encrypt_in: bit_vector5��    (   !                  �                     5�_�   �   �           �   )   "    ����                                                                                                                                                                                                                                                                                                                            [           _           V        f(�0     �   (   *   �      #    signal encrypt_in: bit_vector()5��    (   "                  �                     �    (   &                 �                    �    (   &                 �                    �    (   &                 �                    5�_�   �   �           �   )   /    ����                                                                                                                                                                                                                                                                                                                            [           _           V        f(�5     �   (   *   �      /    signal encrypt_in: bit_vector(511 downto 0)5��    (   /                  �                     5�_�   �   �           �   C   	    ����                                                                                                                                                                                                                                                                                                                            [           _           V        f(�<     �   D   F   �          encrypt_in�   C   F   �              �   C   E   �    5��    C                      l              	       �    C                      l                     �    C                     l              	       �    D                    q                    �    D                 
   q             
       �    D          
          q      
              �    D                 
   q             
       �    D          
       
   q      
       
       �    D          
          q      
              �    D                    q                    5�_�   �   �           �   E       ����                                                                                                                                                                                                                                                                                                                            ]           a           V        f(�E     �   D   F   �              �   D   F   �    5��    D                      m                     �    D                     m                    �    D                    q                    �    D                 	   q             	       �    D          	          q      	              �    D                    q                    �    D                    q                    �    D                    q                    5�_�   �   �           �   E       ����                                                                                                                                                                                                                                                                                                                            ^           b           V        f(�R     �   D   F   �          received_data * 645��    D                     q                     5�_�   �   �           �   F       ����                                                                                                                                                                                                                                                                                                                            ^           b           V        f(�U     �   E   G   �          encrypt_in <= 5��    E                     �                     �    E                    �                    �    E                    �                    �    E                    �                    5�_�   �   �           �   F       ����                                                                                                                                                                                                                                                                                                                            ^           b           V        f(�Z     �   E   G   �          encrypt_in <= received_data5��    E                     �                     5�_�   �   �           �   F       ����                                                                                                                                                                                                                                                                                                                            ^           b           V        f(�c     �   E   G   �          encrypt_in <= 5��    E                     �                     5�_�   �   �           �   F   "    ����                                                                                                                                                                                                                                                                                                                            ^           b           V        f(�o     �   E   G   �      "    encrypt_in <= received_data & 5��    E   "               �  �              �      5�_�   �   �           �   F      ����                                                                                                                                                                                                                                                                                                                            ^           b           V        f(�t     �   E   G   �         encrypt_in <= received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & 5��    E                    �
                     5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            ^           b           V        f(�     �   K   N   �                  msgi =>5��    K                     �
                     �    K                 
   �
             
       �    K          
          �
      
              �    K                    �
                    �    K                                         �    L                                           5�_�   �   �           �   )       ����                                                                                                                                                                                                                                                                                                                            _           c           V        f(݉     �   )   +   �    �   )   *   �    5��    )                      �              1       5�_�   �   �           �   *       ����                                                                                                                                                                                                                                                                                                                            `           d           V        f(݊     �   )   +   �      0    signal encrypt_in: bit_vector(511 downto 0);5��    )                    �                    5�_�   �   �           �   *   #    ����                                                                                                                                                                                                                                                                                                                            `           d           V        f(ݎ     �   )   +   �      1    signal encrypt_out: bit_vector(511 downto 0);5��    )   #                 �                    5�_�   �   �           �   N        ����                                                                                                                                                                                                                                                                                                                            `           d           V        f(ݚ     �   M   P   �       5��    M                      :                     �    M                 
   N             
       �    M          
       
   N      
       
       �    M          
          N      
              �    M                    N                    �    M                    N                    �    M                    N                    �    M                    N                    �    M                     Z                     �    N                      [                     5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                            a           e           V        f(ݪ     �   -   /   �    �   -   .   �    5��    -                      B              $       5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            b           f           V        f(ݯ     �   -   /   �      #    signal finished_receiving: bit;5��    -          	       
   V      	       
       5�_�   �   �           �   P        ����                                                                                                                                                                                                                                                                                                                            b           f           V        f(ݶ    �   O   Q   �       5��    O                      �                     �    O                    �                    �    O                    �                    �    O                    �                    �    O                    �                    5�_�   �   �           �   i   $    ����                                                                                                                                                                                                                                                                                                                            b           f           V        f(��     �   h   j   �      8                        if finished_receiving = '1' then5��    h   $       	          ;      	              �    h                    2                    �    h                    2                    �    h                 
   2             
       �    h          
          2      
              5�_�   �   �           �   p        ����                                                                                                                                                                                                                                                                                                                            o           |           V        f(��     �   n   p   �      8                        if signal_bits_sent < WIDTH then�   o   p          -                            state <= sending;   >                            if signal_bits_sent = WIDTH-1 then   2                                shift_data <= '0';   #                            end if;                           else   .                            state <= stopping;   .                            start_stop <= '1';   #                            -- Data   Q                            parity_bit <= not data_to_parity(word); -- parity bit   2                            parallel_data <= word;   (                            done <= '1';                           end if;    5��    o                            2              �    n           8           �      8               5�_�   �   �           �   n        ����                                                                                                                                                                                                                                                                                                                            n          o           V       f(��     �   m   n          #                    when sending =>    5��    m                      �      %               5�_�   �   �           �   n       ����                                                                                                                                                                                                                                                                                                                            n          n           V       f(��     �   m   o   �      $                    when stopping =>5��    m                    �                    �    m                 
   �             
       �    m          
          �      
              �    m                    �                    �    m                    �                    �    m                    �                    5�_�   �   �           �   j   %    ����                                                                                                                                                                                                                                                                                                                            n          n           V       f(�     �   i   k   �      0                            state <= encrypting;5��    i   %       
          v      
              �    i   %                 v                    �    i   %                 v                    �    i   %                 v                    5�_�   �   �           �   Q        ����                                                                                                                                                                                                                                                                                                                            <          E   
       V   +    f(�     �   Q   S   �    5��    Q                      �              	       �    Q                      �                     5�_�   �   �           �   R        ����                                                                                                                                                                                                                                                                                                                            <          E   
       V   +    f(�     �   R   ]   �    �   R   S   �    5��    R               
       �                    5�_�   �   �           �   S       ����                                                                                                                                                                                                                                                                                                                            <          E   
       V   +    f(�!     �   R   T   �           receiver_component: receiver5��    R                    �                    5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            T          Y          V       f(�k     �   S   U   �              generic map(8)5��    S                     �                     5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            T          Y          V       f(�q     �   S   U   �              generic map(8, 3)5��    S                    �                    5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            T          Y          V       f(�u     �   S   U   �              generic map(8, 10)5��    S                    �                    �    S                    �                    5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            T          Y          V       f(ހ     �   S   U   �              generic map(8, 2)5��    S                      �                      5�_�   �   �           �   V       ����                                                                                                                                                                                                                                                                                                                            T          Y          V       f(ސ     �   U   W   �      "            clock => receiver_clk,5��    U                    4                    �    U                 
   4             
       �    U          
          4      
              �    U                 
   4             
       5�_�   �   �           �   W       ����                                                                                                                                                                                                                                                                                                                            T          Y          V       f(��     �   V   Y   �                  reset,5��    V                    R                     �    W                     _                     �    W                    f                    5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            T          Z          V       f(��     �   .   0   �          �   .   0   �    5��    .                      g                     �    .                     k                     5�_�   �   �           �   f        ����                                                                                                                                                                                                                                                                                                                            U          [          V       f(��     �   f   h   �                      �   f   h   �    5��    f                      �                     �    f                      �                     �    f                    �                    �    f                    �                    �    f                 	   �             	       �    f          	       	   �      	       	       �    f          	          �      	              �    f                    �                    5�_�   �   �           �   g       ����                                                                                                                                                                                                                                                                                                                            U          [          V       f(��     �   f   h   �                      send_data <= 5��    f                     �                     5�_�   �   �           �   g       ����                                                                                                                                                                                                                                                                                                                            U          [          V       f(��     �   f   h   �                      send_data <= ''5��    f                     �                     5�_�   �   �           �   g        ����                                                                                                                                                                                                                                                                                                                            U          [          V       f(��     �   f   h   �                       send_data <= '0'5��    f                      �                     5�_�   �   �           �   y        ����                                                                                                                                                                                                                                                                                                                            U          [          V       f(�     �   y   {   �                                  �   y   {   �    5��    y                                           �    y                                             �    y                 	   +             	       �    y          	       	   +      	       	       �    y          	          +      	              �    y                    +                    5�_�   �   �           �   z   )    ����                                                                                                                                                                                                                                                                                                                            U          [          V       f(�#     �   y   {   �      )                            send_data <= 5��    y   )                  8                     5�_�   �   �           �   z   *    ����                                                                                                                                                                                                                                                                                                                            U          [          V       f(�$     �   y   {   �      +                            send_data <= ''5��    y   *                  9                     5�_�   �   �           �   z   ,    ����                                                                                                                                                                                                                                                                                                                            U          [          V       f(�%     �   y   {   �      ,                            send_data <= '1'5��    y   ,                  ;                     5�_�   �   �           �   Y       ����                                                                                                                                                                                                                                                                                                                            U          [          V       f(�A     �   X   Z   �                  tx_go =>5��    X                     �                     �    X                 	   �             	       �    X          	       	   �      	       	       �    X          	          �      	              �    X                 
   �             
       5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            U          [          V       f(�L     �   Y   [   �      %            serial_data => serial_in,5��    Y                    �                    5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            U          [          V       f(�W     �   /   1   �    �   /   0   �    5��    /                      �              %       5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            V          \          V       f(�Z     �   /   1   �      $    signal finished_encrypting: bit;5��    /          
          �      
              5�_�   �   �           �   [       ����                                                                                                                                                                                                                                                                                                                            V          \          V       f(�e     �   Z   \   �      !            tx_done => serial_in,5��    Z          	          �      	              �    Z                    �                    �    Z                    �                    �    Z                    �                    5�_�   �   �           �   \       ����                                                                                                                                                                                                                                                                                                                            V          \          V       f(�q     �   [   ]   �      '            done => finished_receiving,5��    [                    �                    5�_�   �   �           �   \       ����                                                                                                                                                                                                                                                                                                                            V          \          V       f(�|     �   [   ]   �      '            data => finished_receiving,5��    [                    �                    �    [                    �                    �    [                    �                    �    [                    �                    �    [                    �                    �    [                    �                    5�_�   �   �           �   \       ����                                                                                                                                                                                                                                                                                                                            V          \          V       f(߇     �   [   ]   �                   data => encrypt_out,5��    [                     �                     5�_�   �   �           �   \        ����                                                                                                                                                                                                                                                                                                                            V          \          V       f(߈     �   [   ]   �      "            data => encrypt_out(),5��    [                      �                     �    [   "                 �                    �    [   "                 �                    �    [   "                 �                    5�_�   �   �           �   ]       ����                                                                                                                                                                                                                                                                                                                            V          \          V       f(ߏ     �   \   ]                      data_parity,5��    \                                           5�_�   �   �           �   ]       ����                                                                                                                                                                                                                                                                                                                            V          \          V       f(ߒ     �   \   ^   �      *            parallel_data => received_data5��    \                                        �    \                 	                	       �    \          	                	              �    \                 
                
       �    \                                          5�_�   �   �           �   ]       ����                                                                                                                                                                                                                                                                                                                            V          \          V       f(ߙ     �   \   ^   �      %            serial_o => received_data5��    \                                        �    \                 	                	       �    \          	                	              �    \                 
                
       �    \          
       
         
       
       �    \          
                
              �    \                 
                
       5�_�   �   �           �   ~       ����                                                                                                                                                                                                                                                                                                                            ~          ~   4       v   4    f(߶     �   }      �      \                        if stop_bits_sent < STOP_BITS then -- numero de stop bits arbitrario5��    }                    �                    �    }                    �                    �    }                    �                    �    }                    �                    �    }                    �                    5�_�   �   �           �      %    ����                                                                                                                                                                                                                                                                                                                            ~          ~   4       v   4    f(ߺ     �   ~   �   �      .                            state <= stopping;5��    ~   %                                     5�_�   �   �           �   �   (    ����                                                                                                                                                                                                                                                                                                                            ~          ~   4       v   4    f(��     �      �          .                            start_stop <= '0';5��                                /               5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f(��     �      �                                  else   E                            if start = '1' and serial_data = '0' then   2                                state <= starting;   ,                                done <= '0';       *                                -- Control   4                                start_signal <= '1';   2                                shift_data <= '1';                                else   .                                state <= idle;   ,                                done <= '1';       *                                -- Control   4                                start_signal <= '0';   2                                start_stop <= '0';   2                                shift_data <= '0';5��                                �              5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f(��     �      �          #                            end if;5��                                $               5�_�   �   �   �       �   ~       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f(��     �   }      �    5��    }                      �                     �    }                      �                     5�_�   �   �           �   ~        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f(��     �   }      �                              �   }      �    5��    }                      �                     �    }                      �                     �    }                 	   �             	       �    }          	          �      	              �    }                    �                    5�_�   �   �           �   ~   %    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f(��     �   }      �      %                        send_data <= 5��    }   %                  �                     5�_�   �   �           �   ~   &    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f(��     �   }      �      '                        send_data <= ''5��    }   &                  �                     5�_�   �   �           �   ~   (    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f(��    �   }      �      (                        send_data <= '0'5��    }   (                  �                     5�_�   �   �           �   B       ����                                                                                                                                                                                                                                                                                                                                                             f(�(     �   A   C   �                  reset,5��    A                     \                     �    A                    \                    �    A                    \                    �    A                 	   \             	       5�_�   �   �           �   E       ����                                                                                                                                                                                                                                                                                                                                                             f(�2     �   D   F   �                  data_parity,5��    D                     �                     �    D                 	   �             	       �    D          	       
   �      	       
       �    D          
       
   �      
       
       �    D          
          �      
              �    D                    �                    5�_�   �   �           �   U       ����                                                                                                                                                                                                                                                                                                                                                             f(�H     �   T   V   �          sender_component: receiver5��    T                                        �    T                    !                    5�_�   �   �           �   Y       ����                                                                                                                                                                                                                                                                                                                                                             f(�\    �   X   Z   �                  reset,5��    X                     �                     �    X                    �                    �    X                    �                    �    X                 	   �             	       5�_�   �   �           �   J      ����                                                                                                                                                                                                                                                                                                                                                             f(�y    �   I   K   �         encrypt_in <= received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data5��    I                    A                     5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            L          L          v       f(�     �   K   M   �          encrypt: multisteps�   L   M   �    5��    K          
       
   Q      
       
       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            L          L          v       f(�     �         �          end component�         �          component�         �          �         �    5��                          �                     �                          �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                     	   �             	       �              	          �      	              �                        �                    �                         �                     �                         �                     �                         �                     �                         �                     �                     
   �             
       �              
          �      
              �                     
   �             
       �                        �                     �                         �                    �                         �                    �                         �                     �       
                                       �       	                                        �                        �                    �       
                                       �       	                                        �                     	   �             	       �                                              �                                              �                                              �                                              �                                              �                                              �       
                                       �       	                                        �                     	   �             	       �              	          �      	              �                     
   �             
       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       f(��     �         �    5��                          
                     �                          
                     5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       f(��     �         �    �         �    5��                                        ,       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       f(��     �         �          component multisteps5��              
                
              5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       f(��     �         �    �         �    5��                          �              �       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                       f(��     �         �              clk, rst : in bit;   +        msgi : in bit_vector(511 downto 0);   ,        haso : out bit_vector(255 downto 0);           done : out bit       );�         �      
    port (5��                         �                     �                         
                     �                         )                     �                         Y                     �                         �                     �                         �                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                       f(��     �      *   �    �          �    5��                   
       �              �       5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                       )                 f(��    �       *   �   	           WIDTH: natural := 7;            STOP_BITS : natural := 1       );   	    port(   %        clock, reset, tx_go : in bit;           tx_done : out bit;   /        data : in bit_vector(WIDTH-1 downto 0);           serial_o : out bit       );�      !   �          generic(5��                         �                     �                          �                     �    !                                          �    "                     0                     �    #                     ;                     �    $                     I                     �    %                     s                     �    &                     �                     �    '                     �                     �    (                     �                     5�_�   �              �   O        ����                                                                                                                                                                                                                                                                                                                            O          S           V       f(�     �   M   S          C    receiver_clk <= clock; -- recebe a 5k, mesmo com o clock de 20k       -- receive_clk: slow_clk       --     generic map()   )    --     port map(clock, receiver_clk);    �   S   T   �      C    receiver_clk <= clock; -- recebe a 5k, mesmo com o clock de 20k       -- receive_clk: slow_clk       --     generic map()   )    --     port map(clock, receiver_clk);    �   M   S   �    5��   N              M       `      �       _      �    M                     _                    �    N                     �                    �    O                     �                    �    P                                         5�_�   �                N        ����                                                                                                                                                                                                                                                                                                                            N          R           V       f(�     �   L   R          G        receiver_clk <= clock; -- recebe a 5k, mesmo com o clock de 20k   7                               -- receive_clk: slow_clk   3                               --     generic map()   D                               --     port map(clock, receiver_clk);    �   R   S   �      G        receiver_clk <= clock; -- recebe a 5k, mesmo com o clock de 20k   7                               -- receive_clk: slow_clk   3                               --     generic map()   D                               --     port map(clock, receiver_clk);    �   L   R   �    5��   M              L       _      �       :      5�_�                  M        ����                                                                                                                                                                                                                                                                                                                            M          Q           V       f(�     �   K   Q          G        receiver_clk <= clock; -- recebe a 5k, mesmo com o clock de 20k   7                               -- receive_clk: slow_clk   3                               --     generic map()   D                               --     port map(clock, receiver_clk);    �   Q   R   �      G        receiver_clk <= clock; -- recebe a 5k, mesmo com o clock de 20k   7                               -- receive_clk: slow_clk   3                               --     generic map()   D                               --     port map(clock, receiver_clk);    �   K   Q   �    5��   L              K       :      �             �    K                                         �    L                     R                    �    M                     �                    �    N                     �                    5�_�                 L        ����                                                                                                                                                                                                                                                                                                                            L          P           V       f(�     �   J   P          C    receiver_clk <= clock; -- recebe a 5k, mesmo com o clock de 20k   3                           -- receive_clk: slow_clk   /                           --     generic map()   @                           --     port map(clock, receiver_clk);    �   P   Q   �      C    receiver_clk <= clock; -- recebe a 5k, mesmo com o clock de 20k   3                           -- receive_clk: slow_clk   /                           --     generic map()   @                           --     port map(clock, receiver_clk);    �   J   P   �    5��   K              J             �       �      5�_�                 K        ����                                                                                                                                                                                                                                                                                                                            K          O           V       f(�     �   I   O          C    receiver_clk <= clock; -- recebe a 5k, mesmo com o clock de 20k   3                           -- receive_clk: slow_clk   /                           --     generic map()   @                           --     port map(clock, receiver_clk);    �   O   P   �      C    receiver_clk <= clock; -- recebe a 5k, mesmo com o clock de 20k   3                           -- receive_clk: slow_clk   /                           --     generic map()   @                           --     port map(clock, receiver_clk);    �   I   O   �    5��   J              I       �      �       �      5�_�               K       ����                                                                                                                                                                                                                                                                                                                            K          M                 f(��     �   J   L   �      3                           -- receive_clk: slow_clk5��    J                                          5�_�                 L       ����                                                                                                                                                                                                                                                                                                                            K          M                 f(��     �   K   M   �      /                           --     generic map()5��    K                     7                     5�_�                 M       ����                                                                                                                                                                                                                                                                                                                            K          M                 f(��   	 �   L   N   �      @                           --     port map(clock, receiver_clk);5��    L                     P                     5�_�    	             J       ����                                                                                                                                                                                                                                                                                                                            K          M                 f(��     �   I   K   �      C    receiver_clk <= clock; -- recebe a 5k, mesmo com o clock de 20k5��    I                     �      D       G       5�_�    
          	   M       ����                                                                                                                                                                                                                                                                                                                            K          M          V       f(��     �   J   N   �          -- receive_clk: slow_clk       --     generic map()   )    --     port map(clock, receiver_clk);5��    J                           `       W       5�_�  	            
   K       ����                                                                                                                                                                                                                                                                                                                            K          M          V       f(��     �   J   L   �          receive_clk: slow_clk5��    J                     2                     5�_�  
               L       ����                                                                                                                                                                                                                                                                                                                            K          M          V       f(��     �   K   M   �              generic map()5��    K                  %   I              %       5�_�                 L   :    ����                                                                                                                                                                                                                                                                                                                            K          M          V       f(�>     �   K   M   �      :        generic map()   -- Converte clock de 50M pra 192005��    K   :                  n                     5�_�                 L       ����                                                                                                                                                                                                                                                                                                                            K          M          V       f(�B     �   K   M   �      <        generic map()   -- Converte clock de 50M pra 19200Hz5��    K                     H                     5�_�                 O       ����                                                                                                                                                                                                                                                                                                                            K          M          V       f(�i     �   N   O              -- Clocks do judge5��    N                      �                     5�_�                 J       ����                                                                                                                                                                                                                                                                                                                            K          M          V       f(�k     �   I   K   �    �   J   K   �    5��    I                      �                     5�_�                 J       ����                                                                                                                                                                                                                                                                                                                            L          N          V       f(�m     �   I   K   �          -- Clocks do judge5��    I                     �                     5�_�                 Q   +    ����                                                                                                                                                                                                                                                                                                                            L          N          V       f(�u     �   P   R   �      +        generic map(2) -- clock divido em 45��    P   +                                       �    P   *                                     �    P   1                                     �    P   1                                     �    P   1              
                
       �    P   :                                     �    P   <                 !                    5�_�                 Q       ����                                                                                                                                                                                                                                                                                                                            L          N          V       f(�     �   P   R   �      H        generic map(2) -- clock divido em 2 para judge e 5208 para placa5��    P                    �                    �    P                    �                    �    P                    �                    �    P                    �                    5�_�                 K   F    ����                                                                                                                                                                                                                                                                                                                            L          N          V       f(�     �   J   L   �      F    -- receiver_clk <= clock; -- recebe a 5k, mesmo com o clock de 20k5��    J   !       %                %              5�_�                 M   @    ����                                                                                                                                                                                                                                                                                                                            L          N          V       f(�   
 �   L   N   �      @        generic map(1302)   -- Converte clock de 50M pra 19200Hz5��    L   @                  �                     5�_�                 {       ����                                                                                                                                                                                                                                                                                                                            L          N          V       f(��    �   z   {          "                serial_out <= '1';5��    z                      [      #               5�_�                 D       ����                                                                                                                                                                                                                                                                                                                            E          E          V       f(�     �   C   E   �    �   D   E   �    5��    C                      d              %       5�_�                 D       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(�     �   C   E   �      $    signal finished_encrypting: bit;5��    C                    o                    5�_�                 }       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(�     �   }      �                      �   }      �    5��    }                      �                     �    }                     �                     �    }                     �                     �    }                     �                     �    }                     �                     �    }                    �                    �    }                    �                    �    }                    �                    5�_�                 ~   $    ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(�     �   }      �      $                start_encrypting <= 5��    }   $                  �                     5�_�                 ~   %    ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(�     �   }      �      &                start_encrypting <= ''5��    }   %                  �                     5�_�                 ~   '    ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(�     �   }      �      '                start_encrypting <= '0'5��    }   '                  �                     5�_�                 �   '    ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   �   �   �    �   �   �   �    5��    �                      �              )       5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   �   �   �    5��    �                      �                     �    �                     �                    �    �                      �                     5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   �   �   �      (                start_encrypting <= '0';5��    �                     
                     5�_�                  �       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   �   �          4                            start_encrypting <= '0';5��    �                      �      5               5�_�    !              �        ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   �   �   �    �   �   �   �    5��    �                      z              5       5�_�     "          !   �       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   �   �   �      4                            start_encrypting <= '0';5��    �                     �                     5�_�  !  #          "   �       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   �   �          0                        start_encrypting <= '0';5��    �                      z      1               5�_�  "  $          #   �        ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   �   �   �    �   �   �   �    5��    �                      �              1       5�_�  #  %          $   �       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   �   �   �      0                        start_encrypting <= '0';5��    �                     �                     5�_�  $  &          %   �       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   �   �   �    5��    �                      +                     �    �                      +                     5�_�  %  '          &   �        ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   �   �   �    �   �   �   �    5��    �                      ,              1       5�_�  &  (          '   �       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   �   �   �      0                        start_encrypting <= '0';5��    �                     D                     5�_�  '  )          (   �        ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   �   �           5��    �                      +                     5�_�  (  *          )   �   1    ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   �   �   �      4                            start_encrypting <= '0';5��    �   1                 \                    5�_�  )  +          *   �   1    ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(�,     �   �   �          4                            start_encrypting <= '0';5��    �                            5               5�_�  *  ,          +   �   )    ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(�/     �   �   �   �    �   �   �   �    5��    �                      .              5       5�_�  +  -          ,   �        ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(�1     �   �   �           5��    �                      c                     5�_�  ,  .          -   f       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(�E     �   e   g   �                  reset,5��    e                     '                     �    e                     -                     �    e                     ,                     �    e                    +                    �    e                    +                    �    e                    +                    5�_�  -  /          .   f       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(�M     �   e   g   �      &            reset => start_encrypting,5��    e                    "                    �    e                     #                     �    e                    "                    �    e                    "                    �    e                    "                    5�_�  .  7          /   f       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(�T    �   e   g   �      $            rst => start_encrypting,5��    e                     )                     5�_�  /  8  0      7   B       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f)}     �   B   D   �          �   B   D   �    5��    B                      @                     �    B                     D                     5�_�  7  9          8   C       ����                                                                                                                                                                                                                                                                                                                            G          G          V       f)�     �   B   C              signal done5��    B                      @                     5�_�  8  :          9   D       ����                                                                                                                                                                                                                                                                                                                            F          F          V       f)�     �   C   E   �    5��    C                      d                     �    C                      d                     5�_�  9  ;          :   F       ����                                                                                                                                                                                                                                                                                                                            G          G          V       f)�     �   E   F          $    signal finished_encrypting: bit;5��    E                      �      %               5�_�  :  <          ;   D        ����                                                                                                                                                                                                                                                                                                                            F          F          V       f)�     �   C   E   �    �   D   E   �    5��    C                      d              %       5�_�  ;  =          <   H       ����                                                                                                                                                                                                                                                                                                                            G          G          V       f)�     �   G   H          !    signal finished_sending: bit;5��    G                      �      "               5�_�  <  >          =   E        ����                                                                                                                                                                                                                                                                                                                            G          G          V       f)�     �   D   F   �    �   E   F   �    5��    D                      �              "       5�_�  =  @          >   C       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)�     �   B   D   �          signal _receiving: bit;�   B   F   �      #    signal finished_receiving: bit;   $    signal finished_encrypting: bit;   !    signal finished_sending: bit;5��    B                     K                     �    C                     g                     �    D                     �                     �    B                     K                     �    C                     k                     �    D                     �                     5�_�  >  A  ?      @   \        ����                                                                                                                                                                                                                                                                                                                            E          C                 f)�     �   �   �          R                        if finished_sending then -- numero de stop bits arbitrario�   �   �          9                        if finished_encrypting = '1' then�   �   �          8                        if finished_receiving = '1' then�   r   t          (            tx_done => finished_sending,�   i   k          '            done => finished_encrypting�   [   ]   �      '            done => finished_receiving,5��    [                    0	                    �    i                    �                    �    r                    ~                    �    �                    �                    �    �                    �                    �    �                    �                    5�_�  @  B          A   H       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)�     �   G   I   �          signal send_data: bit;5��    G                     �                     5�_�  A  C          B   H       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)�     �   G   I   �          signal send: bit;5��    G                     �                     5�_�  B  D          C   H       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)�     �   G   I   �          signal start_send: bit;5��    G                     �                     5�_�  C  E          D   r       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)�     �   q   s   �                  tx_go => send_data,5��    q          	          `      	              �    q                     b                     �    q                     a                     �    q                    `                    �    q                    `                    �    q                    `                    5�_�  D  F          E   ~       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)�     �   }      �      !                send_data <= '0';5��    }          	          �      	              �    }                     �                     �    }                     �                     �    }                    �                    �    }                    �                    �    }                    �                    5�_�  E  G          F   �       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)�     �   �   �   �      -                            send_data <= '1';5��    �          	          1      	              �    �                     3                     �    �                     2                     �    �                    1                    �    �                    1                    �    �                    1                    �    �                    1                    5�_�  F  J          G   �       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)�    �   �   �   �      )                        send_data <= '0';5��    �          	          �      	              �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�  G  K  H      J   �       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)�     �   �   �          4                            start_encrypting <= '0';5��    �                      5      5               5�_�  J  L          K   �       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)�    �   �   �   �    �   �   �   �    5��    �                      G              5       5�_�  K  M          L   �       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)"     �   �   �          4                            start_encrypting <= '0';5��    �                      G      5               5�_�  L  N          M   �       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)"    �   �   �   �    �   �   �   �    5��    �                      5              5       5�_�  M  O          N   �       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)#�     �   �   �          -                        start_sending <= '0';5��    �                      �      .               5�_�  N  P          O   �        ����                                                                                                                                                                                                                                                                                                                            E          C                 f)#�     �   �   �   �    �   �   �   �    5��    �                      <              .       5�_�  O  Q          P   �       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)#�     �   �   �   �      -                        start_sending <= '0';5��    �                     T                     5�_�  P              Q   �        ����                                                                                                                                                                                                                                                                                                                            E          C                 f)#�    �   �   �           5��    �                      �                     5�_�  G  I      J  H   �       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)�     �   �   �        5��    �                      5      5               5�_�  H              I   �       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)�     �   �   �   �    �   �   �   �      4                            start_encrypting <= '0';5��    �                      G              5       5�_�  >          @  ?   C       ����                                                                                                                                                                                                                                                                                                                            E          C                 f)�     �   B   D   �          signal don_receiving: bit;5��    B                     N                     5�_�  /  1      7  0   Z        ����                                                                                                                                                                                                                                                                                                                            F          F          V       f(��     �   Y   Z   �                  �   Y   [   �                  start =>5��    Y                      	                     �    Y                     	                     �    Y                    	                    5�_�  0  2          1   C       ����                                                                                                                                                                                                                                                                                                                            G          G          V       f(��     �   C   D   �    �   B   C   �      !    signal start_encrypting: bit;5��    B                      @              "       5�_�  1  3          2   C       ����                                                                                                                                                                                                                                                                                                                            G          G          V       f(��     �   B   D   �           signal start_receiving: bit;5��    B          
          Q      
              �    B                     X                     �    B                    W                    5�_�  2  4          3   [       ����                                                                                                                                                                                                                                                                                                                            G          G          V       f(��     �   Z   \   �      %            start => start_receiving,5��    Z                     6	                     �    Z                     :	                     �    Z                     9	                     �    Z                     8	                     �    Z                    7	                    �    Z   #                  E	                     �    Z   "                  D	                     �    Z   !                  C	                     �    Z                      B	                     �    Z                     A	                     �    Z                     @	                     �    Z                     ?	                     �    Z                     >	                     �    Z                     =	                     �    Z                     <	                     �    Z                     ;	                     �    Z                     :	                     �    Z                     9	                     �    Z                     8	                     �    Z                    7	                    �    Z                    7	                    �    Z                    7	                    5�_�  3  5          4          ����                                                                                                                                                                                                                                                                                                                            G          G          V       f(�    �         �      5            clock, reset, start, serial_data: in bit;5��                         F                     5�_�  4  6          5   �       ����                                                                                                                                                                                                                                                                                                                            G          G          V       f(�(     �   �   �   �    �   �   �   �      (                start_encrypting <= '0';5��    �                      -              )       5�_�  5              6   �       ����                                                                                                                                                                                                                                                                                                                            G          G          V       f(�,     �   �   �   �      '                start_receiving <= '0';5��    �          	           D      	               �    �                    C                    �    �                     F                     �    �                     E                     �    �                     D                     �    �                     C                     �    �                     B                     �    �                     A                     �    �                     @                     �    �                     ?                     �    �                     >                     �    �                    =                    �    �                    =                    �    �                    =                    5�_�                 K       ����                                                                                                                                                                                                                                                                                                                            J          N           V       f(��     �   J   L   �               -- receive_clk: slow_clk5��    J                                          5�_�   �       �   �   �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f(��     �   �   �   �                              �   �   �   �                              se5��    �                      4                     �    �                     L                     5�_�   �           �   �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f(��     �      �   �                                  �      �   �           5��                                               �                                             �                                               �                                              �    �                                           5�_�   �           �   �   W        ����                                                                                                                                                                                                                                                                                                                            S           W           V        f(�k     �   W   X   �    �   W   X   �      %                    when receiving =>   8                        if finished_receiving = '1' then   0                            state <= encrypting;                               end if;5��    W                      w              �       5�_�   �           �   �   Y       ����                                                                                                                                                                                                                                                                                                                            O   !       R          V   !    f(�     �   X   [        5��    X                      k      W               5�_�   M           O   N          ����                                                                                                                                                                                                                                                                                                                                         #       V   #    f(�r     �          m          _clk: sender_clk5��                                              5�_�   =           ?   >          ����                                                                                                                                                                                                                                                                                                                                                             f(��     �         V    �         V      #    signal receiversender_clk: bit;5��                         �                      5�_�             !             ����                                                                                                                                                                                                                                                                                                                                                             f'ז     �                        serial_ i n : in b i t ;5��                         M                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'ח     �                       serial_  n : in b i t ;5��                         O                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f'ח     �                       serial_   : in b i t ;5��                         P                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f'ח     �                       serial_    in b i t ;5��                         Q                      5�_�                             ����                                                                                                                                                                                                                                                                                                                                                             f'ח     �                       serial_    n b i t ;5��                         R                      5�_�                          ����                                                                                                                                                                                                                                                                                                                                                             f'ׁ     �                ent  t y sha256_1b i s5��                                                5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f'ׂ     �                ent   y sha256_1b i s5��                                                5��