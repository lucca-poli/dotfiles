Vim�UnDo� �Y]���]��1�
�`�3٫�M�*_vZ��?��   i                                   f(AI    _�                     B        ����                                                                                                                                                                                                                                                                                                                                                             f�x    �   B            �   B            5��    B                      �              $      5�_�                   D       ����                                                                                                                                                                                                                                                                                                                                                             f�     �   C   E   `      "use IEEE.NUMERIC_BIT_UNSIGNED.ALL;5��    C          	           �      	               5�_�                    S       ����                                                                                                                                                                                                                                                                                                                                                             f�    �   R   T   `      "use IEEE.NUMERIC_BIT_UNSIGNED.ALL;5��    R          	           �      	               5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f>*    �          `    �         `    5��                                                 5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             fI     �      
          %architecture behavioral of somador is�                end entity somador;�          t      entity somador is5��                                              �                        �                     �                        �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             fI     �         t      '        A : in bit_vector(31 downto 0);5��                        %                     5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                             fI     �         t      '        B : in bit_vector(31 downto 0);5��                        M                     5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                             fI	     �         t      '        S : out bit_vector(31 downto 0)5��                        u                     5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                             fI     �         t      +        S(i) <= A(i) xor B(i) xor carry(i);5��                        4                    5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                             fI    �         t      +    S(31) <= A(31) xor B(31) xor carry(31);5��                        �                    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f�J     �      
          %architecture behavioral of adder32 is�                end entity adder32;�          t      entity adder32 is5��                      	                 	       �                     	   �              	       �                     	   �              	       5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        f�P    �                 entity somador32 is   
    port (   '        a : in bit_vector(31 downto 0);   '        b : in bit_vector(31 downto 0);   '        r : out bit_vector(31 downto 0)       );   end entity somador32;       'architecture behavioral of somador32 is   +    signal carry : bit_vector(31 downto 0);   begin   "    sum: for i in 0 to 30 generate   +        r(i) <= A(i) xor B(i) xor carry(i);   T        carry(i+1) <= (A(i) and B(i)) or (A(i) and carry(i)) or (B(i) and carry(i));       end generate;       +    r(31) <= A(31) xor B(31) xor carry(31);          end architecture behavioral;    5��                                                 5�_�                    
        ����                                                                                                                                                                                                                                                                                                                                       `           V        f��     �   
   k   `    �   
      `    5��    
               `       �               �      5�_�                            ����                                                                                                                                                                                                                                                                                                                                       �           V        f�w     �              �   library ieee;   use ieee.numeric_bit.all;       entity ch is   	port (   )    	x, y, z: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end ch;       library ieee;   use ieee.numeric_bit.all;       entity ch is   	port (   )    	x, y, z: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end ch;       architecture arch1 of ch is   0	signal op1, op2, op3 : bit_vector(31 downto 0);   begin   	op1 <= x and y;       op2 <= (not x) and z;       op3 <= op1 xor op2;        q <= op3;   
end arch1;       entity maj is   	port (   )    	x, y, z: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end maj;       architecture arch2 of maj is   4	signal op1, op2, op3, op4: bit_vector(31 downto 0);   begin   	op1 <= x and y;       op2 <= x and z;       op3 <= y and z;        op4 <= op1 xor op2 xor op3;        q <= op4;   
end arch2;       library ieee;   use ieee.numeric_bit.all;       entity sum0 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   	end sum0;       architecture arch3 of sum0 is   begin   1    q <= (x ror 2) xor (x ror 13) xor (x ror 22);   
end arch3;       library ieee;   use ieee.numeric_bit.all;       entity sum1 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   	end sum1;       architecture arch4 of sum1 is   begin   1    q <= (x ror 6) xor (x ror 11) xor (x ror 25);   
end arch4;       library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity sigma0 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end sigma0;       architecture arch5 of sigma0 is   begin   0    q <= (x ror 7) xor (x ror 18) xor (x srl 3);   
end arch5;       library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity sigma1 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end sigma1;       architecture arch6 of sigma1 is   begin   2    q <= (x ror 17) xor (x ror 19) xor (x srl 10);   
end arch6;       architecture arch1 of ch is   0	signal op1, op2, op3 : bit_vector(31 downto 0);   begin   	op1 <= x and y;       op2 <= (not x) and z;       op3 <= op1 xor op2;        q <= op3;   
end arch1;       entity maj is   	port (   )    	x, y, z: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end maj;       architecture arch2 of maj is   4	signal op1, op2, op3, op4: bit_vector(31 downto 0);   begin   	op1 <= x and y;       op2 <= x and z;       op3 <= y and z;        op4 <= op1 xor op2 xor op3;        q <= op4;   
end arch2;       library ieee;   use ieee.numeric_bit.all;       entity sum0 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   	end sum0;       architecture arch3 of sum0 is   begin   1    q <= (x ror 2) xor (x ror 13) xor (x ror 22);   
end arch3;       library ieee;   use ieee.numeric_bit.all;       entity sum1 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   	end sum1;       architecture arch4 of sum1 is   begin   1    q <= (x ror 6) xor (x ror 11) xor (x ror 25);   
end arch4;       library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity sigma0 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end sigma0;       architecture arch5 of sigma0 is   begin   0    q <= (x ror 7) xor (x ror 18) xor (x srl 3);   
end arch5;       library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity sigma1 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end sigma1;       architecture arch6 of sigma1 is   begin   2    q <= (x ror 17) xor (x ror 19) xor (x srl 10);   
end arch6;    5��            �                      h             5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        f�y     �                   �               5��                    a                       �      5�_�                    b        ����                                                                                                                                                                                                                                                                                                                                                  V        f�z     �   a   b           5��    a                      �                     5�_�                    a        ����                                                                                                                                                                                                                                                                                                                                                  V        f�{    �   `   a           5��    `                      �                     5�_�                    F        ����                                                                                                                                                                                                                                                                                                                            F          `           V       f�n     �   E   F          entity sigma0 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end sigma0;       architecture arch5 of sigma0 is   begin   0    q <= (x ror 7) xor (x ror 18) xor (x srl 3);   
end arch5;       library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity sigma1 is   	port (   #    	x: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)   
        );   end sigma1;       architecture arch6 of sigma1 is   begin   2    q <= (x ror 17) xor (x ror 19) xor (x srl 10);   
end arch6;    5��    E                      �      �              5�_�                    C        ����                                                                                                                                                                                                                                                                                                                            F          F           V       f�o    �   B   C          library IEEE;   use IEEE.NUMERIC_BIT.ALL;    5��    B                      �      )               5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f(A6     �          B    5��                                                  5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f(AF     �       (   D       �         D    �          C    5��                                                  �                    &                       �      5�_�                     '        ����                                                                                                                                                                                                                                                                                                                                                             f(AH    �   &   '           5��    &                      �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f(A;     �          C       �         D    �          D      Hhttps://drive.google.com/drive/folders/1Rg1G8QwLyDoD_2JOD1SH4AR_5yNKS2pi5��                                                  �                        H                   H       5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f(A8     �         C    �          C       5��                                                  5�_�                    D       ����                                                                                                                                                                                                                                                                                                                                                             f�
     �   C   E   `      use IEEE.NUMERIC_BITALL;5��    C          
           �      
               5��