Vim�UnDo� ���:����@�Q�	I�7��LS>�nlj���   G           /                       e�=K    _�                            ����                                                                                                                                                                                                                                                                                                                                                             e�9�     �                   �               5��                   G                      �      5�_�                       	    ����                                                                                                                                                                                                                                                                                                                                                             e�9�     �         H          dut: ch5��       	                 �                    5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                             e�9�     �   	      H          component ch5��    	                    �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�9�     �         H      entity ch_tb is end;5��                        E                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�9�    �      	   H      architecture dut of ch_tb is5��                        i                     �                         k                      �                         j                      �                        i                     �                         k                      �                         j                      �                        i                     �                        i                     �                        i                     �                        i                     5�_�                       /    ����                                                                                                                                                                                                                                                                                                                            7          7          v       e�<�    �         H      =        file tb_file : text open read_mode is "cases_ch.dat";5��       /                 �                    5�_�                             ����                                                                                                                                                                                                                                                                                                                                                  V   ;    e�=J    �                  5��                                                  5�_�                             ����                                                                                                                                                                                                                                                                                                                                                             e�9�     �              �                     use ieee.numeric_bit.ALL;5��                                                5��