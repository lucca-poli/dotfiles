Vim�UnDo� z^��J�T7+��tMl�v!�䇰iG1E�   �   +                        if start = '1' then   �   &                       f�     _�                    8        ����                                                                                                                                                                                                                                                                                                                                                             fMl     �   9   G   �       �   :   ;   �    �   8   ;   �       �   8   :   �    5��    8                      (                     �    8                      (                     �    9                     )              �      5�_�                    0       ����                                                                                                                                                                                                                                                                                                                                                             fMw     �   /   1   �               STOP_BITS : natural := 15��    /          	          [      	              �    /                 	   [             	       �    /          	       	   [      	       	       �    /          	          [      	              �    /                 	   [             	       5�_�                    0       ����                                                                                                                                                                                                                                                                                                                                                             fM     �   /   1   �               CLOCK_MUL : natural := 15��    /                     d                     5�_�                    /       ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   .   0   �              PARITY : natural := 1;5��    .                     B                     5�_�                    -       ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   ,   .   �      #        POLARITY : boolean := TRUE;5��    ,                                          5�_�                    0       ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   /   1   �              CLOCK_MUL: natural := 15��    /                    o                    5�_�      	              3       ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   2   4   �      %        clock, reset, tx_go : in bit;5��    2                    �                    5�_�      
           	   3   (    ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   2   4   �      2        clock, reset, start, serial_data : in bit;5��    2   (                  �                     5�_�   	              
   4       ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   3   5   �              tx_done : out bit;5��    3                 	   �             	       �    3                 
   �             
       5�_�   
                 4       ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   3   5   �      #        done, parity_bit : out bit;5��    3                     �                     5�_�                    5       ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   4   6   �      /        data : in bit_vector(WIDTH-1 downto 0);5��    4                    �                    �    4                 
   �             
       5�_�                    5       ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   4   6   �      8        parallel_data : in bit_vector(WIDTH-1 downto 0);5��    4                    �                    5�_�                    5       ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   4   6   �      9        parallel_data : out bit_vector(WIDTH-1 downto 0);5��    4                     �                     5�_�                    6       ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   5   6                  serial_o : out bit5��    5                                           5�_�                    7       ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   6   8   �      end serial_out;5��    6                    "                    5�_�                    +       ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   *   ,   �      entity serial_out is5��    *                    �                    5�_�                    7       ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   6   8   �      end serial_in;5��    6          	                	              �    6                                          �    6                                        5�_�                    9        ����                                                                                                                                                                                                                                                                                                                                                             fM�     �   8   9          !e n t i t y s e r i a l _ i n i s   g en e r ic (   POLARITY : boolean := TRUE;   WIDTH: n a t u r a l := 8 ;   PARITY : n a t u r a l := 1 ;   CLOCK_MUL: p o s i t i v e := 4   ) ;   po r t (   Bclock , r e s e t , s t a r t , s e r i a l _ d a t a : in b i t ;   (done , p a r i t y _ b i t : out b i t ;   Hp a r a l l e l _ d a t a : out b i t _ v e c t o r (WIDTH−1 downto 0)   ) ;   end s e r i a l _ i n ;    5��    8                      #      �              5�_�                    9       ����                                                                                                                                                                                                                                                                                                                                                             fM�    �   8   :   �      (architecture Behavioral of serial_out is5��    8          
          >      
              �    8                     @                     �    8                     ?                     �    8                 	   >             	       �    8          	       	   >      	       	       �    8          	          >      	              �    8                 	   >             	       5�_�                    F        ����                                                                                                                                                                                                                                                                                                                                                             fPa     �   E   F       	   M    function data_to_parity(data: bit_vector(WIDTH-1 downto 0)) return bit is   ,        variable xor_result: bit := data(0);   	begin   "        for i in 1 to WIDTH-1 loop   1            xor_result := xor_result xor data(i);           end loop;           return xor_result;   	end function;    5��    E       	               �                    5�_�                    I        ����                                                                                                                                                                                                                                                                                                                                                             fPw     �   I   K   �          �   I   K   �    5��    I                      =                     �    I                     A                     �    I                     P                     �    I                    O                    �    I                    [                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             fQi     �          �    5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             fQk     �          �       �         �    �          �    5��                                                  �                                           O      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             fQm     �                 5��                          O                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             fQw     �          �      entity shift_reg512 is5��                                              5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             fQ}     �      	   �      end entity shift_reg512;5��                        �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             fQ     �      	   �      end entity shift_reg8;5��              
           �       
               5�_�                       
    ����                                                                                                                                                                                                                                                                                                                                                             fQ�     �      	   �      end entity ;5��       
                  �                      5�_�                    
   "    ����                                                                                                                                                                                                                                                                                                                                                             fQ�     �   	      �      (architecture Behavior of shift_reg512 is5��    	   "                 �                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             fQ�     �   
      �      ,   signal vector: bit_vector(511 downto 0); 5��    
                                        5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                                             fQ�     �         �      '        d: in bit_vector(511 downto 0);5��                        �                     5�_�       "           !          ����                                                                                                                                                                                                                                                                                                                                                             fQ�     �         �      '        q: out bit_vector(511 downto 0)5��                        �                     5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                                                             fQ�     �         �      )        data: in bit_vector(31 downto 0);5��                        ^                     5�_�   "   $           #          ����                                                                                                                                                                                                                                                                                                                                                             fQ�     �                (        data: in bit_vector(7 downto 0);5��                          B       )               5�_�   #   %           $      	    ����                                                                                                                                                                                                                                                                                                                                                             fR    �                
    port (   !        rst, clk, enable: in bit;5��                                               5�_�   $   &           %          ����                                                                                                                                                                                                                                                                                                                                                             f�8     �         �          rst, clk, enable: in bit;5��                         $                      5�_�   %   '           &          ����                                                                                                                                                                                                                                                                                                                                                             f�:     �         �          �         �    5��                          B               	       �                         B                     �                     	   N              	       5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �         �      2            vector <= vector(479 downto 0) & data;5��                        �                    �                         �                     �                        �                    �       !                  �                     �                          �                     �                         �                     �                         �                     �                        �                    �       "                  �                     �       !                  �                     �                          �                     �                         �                     �                         �                     �                        �                    5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �         �      0            vector <= vector(6 downto 0) & data;5��                        �                    5�_�   (   *           )      &    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �         �      0            vector <= vector(7 downto 0) & data;5��       &                 �                    5�_�   )   +           *      (    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �         �      0            vector <= vector(7 downto 1) & data;5��       (                  �                     5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �         �      )            vector <= vector(7 downto 1);5��                         �                     5�_�   +   -           ,   d   -    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f�     �   c   e   �      .    signal word: bit_vector(WIDTH-1 downto 0);5��    c   -                  ^	                     �    c   1                  b	                     5�_�   ,   .           -   d   1    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f�     �   c   e   �      2    signal word: bit_vector(WIDTH-1 downto 0) := ;5��    c   1                  b	                     5�_�   -   /           .   d   2    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f�     �   c   e   �      4    signal word: bit_vector(WIDTH-1 downto 0) := ();5��    c   2                  c	                     �    c   2                 c	                    �    c   2                 c	                    �    c   2                 c	                    �    c   2                 c	                    5�_�   .   0           /          ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f�@     �         �                  vector <= d;5��                         f                     5�_�   /   1           0          ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f�A     �         �                  vector <= ;5��                         f                     5�_�   0   2           1          ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f�A     �         �                  vector <= ();5��                         g                     �                        g                    �                        g                    �                        g                    �                        g                    5�_�   1   3           2   P   8    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f�T     �   O   Q   �      8        parallel_data: out bit_vector(WIDTH-1 downto 0);5��    O   7                  >                     5�_�   2   4           3   r       ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �   q   s   �      8        generic map(STOP_BITS+1) -- Stop bits and parity5��    q          	          �
      	              5�_�   3   5           4   s       ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f�p     �   u   w   �              port�   t   w   �          incoming_data: shift_reg8�   s   v   �              �   s   u   �    5��    s                      ^              	       �    s                      ^                     �    s                     ^              	       �    t                    c                    �    t                     o                     �    t                    n                    �    t                     t                     �    t                     s                     �    t                 
   r             
       �    t          
          r      
              �    t                 
   r             
       �    t                    |                     �    u                     �                     �    u   	                 �                    �    u                    �                    �    u                    �                    �    u                    �                    5�_�   4   6           5   v       ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �   u   w   �              port map5��    u                     �                     5�_�   5   7           6          ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �                %        d: in bit_vector(7 downto 0);5��                          X       &               5�_�   6   8           7   
   (    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �   	      �      *   signal vector: bit_vector(7 downto 0); 5��    	   (                  �                      5�_�   7   9           8   
   ,    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �   	      �      .   signal vector: bit_vector(7 downto 0) := ; 5��    	   ,                  �                      5�_�   8   :           9   
   -    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �   	      �      0   signal vector: bit_vector(7 downto 0) := (); 5��    	   -                  �                      �    	   -                 �                     �    	   -                 �                     �    	   -                 �                     �    	   -                 �                     5�_�   9   ;           :   u       ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �   t   v   �              port map()5��    t                     {                     �    t                    {                    �    t                    {                    �    t                 
   {             
       �    t                    �                    �    t                    �                    �    t                 
   �             
       5�_�   :   <           ;   u   "    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �   t   v   �      #        port map(reset, clock, en,)5��    t   "                  �                     5�_�   ;   =           <   u   )    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �   t   v   �      *        port map(reset, clock, en, data, )5��    t   )                  �                     5�_�   <   >           =   c   -    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �   b   d   �      A    signal word: bit_vector(WIDTH-1 downto 0) := (others => '0');5��    b   -                  X	                     5�_�   =   ?           >   h   -    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �   h   j   �          �   h   j   �    5��    h                      
                     �    h                  
   
              
       �    h                     
                     �    h                    
                    5�_�   >   @           ?   i       ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f��     �   h   j   �          signal shift_data: bit;5��    h                     !
                     �    h                     !
                     5�_�   ?   A           @   v       ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f�     �   u   w   �      .        port map(reset, clock, en, data, word)5��    u                    �                    �    u                 
   �             
       �    u          
       
   �      
       
       �    u          
       
   �      
       
       �    u          
          �      
              �    u                 
   �             
       5�_�   @   B           A   v   +    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f�     �   u   w   �      6        port map(reset, clock, shift_data, data, word)5��    u   +                 �                    �    u   +                 �                    �    u   +              	   �             	       �    u   +       	       	   �      	       	       �    u   +       	          �      	              �    u   +              	   �             	       5�_�   A   C           B   v   +    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f�     �   u   w   �      ;        port map(reset, clock, shift_data, serial_in, word)5��    u   +       	          �      	              �    u   ,                 �                    �    u   +                 �                    �    u   +                 �                    �    u   +                 �                    �    u   +                 �                    5�_�   B   D           C   v   =    ����                                                                                                                                                                                                                                                                                                                                         +       v   +    f�%    �   u   w   �      =        port map(reset, clock, shift_data, serial_data, word)5��    u   =                  �                     5�_�   C   E           D   �       ����                                                                                                                                                                                                                                                                                                                                                             f�e     �   �   �   �      +                        if tx_go = '1' then5��    �                    ~                    �    �                     �                     �    �                                          �    �                    ~                    �    �                    ~                    �    �                    ~                    �    �   "                  �                     �    �   !                  �                     �    �                      �                     5�_�   D   F           E   �       ����                                                                                                                                                                                                                                                                                                                                                             f�     �   �   �   �      +                            tx_done <= '0';5��    �                    �                    5�_�   E   G           F   �       ����                                                                                                                                                                                                                                                                                                                                                             f�>     �   �   �          (                word <= (others => '0');5��    �                      �      )               5�_�   F   H           G   }       ����                                                                                                                                                                                                                                                                                                                                                             f�Q     �   |   ~   �                      tx_done <= '1';5��    |                     T                     5�_�   G   I           H   }       ����                                                                                                                                                                                                                                                                                                                                                             f�R     �   |   ~   �                      x_done <= '1';5��    |                     T                     5�_�   H   J           I   }       ����                                                                                                                                                                                                                                                                                                                                                             f�R     �   |   ~   �                      _done <= '1';5��    |                     T                     5�_�   I   K           J   ~       ����                                                                                                                                                                                                                                                                                                                                                             f�S     �   }      �                       serial_o <= '1';5��    }                    q                    �    }                     u                     �    }                     t                     �    }                     s                     �    }                     r                     �    }                    q                    �    }                     v                     �    }                     u                     �    }                     t                     �    }                     s                     �    }                     r                     �    }                 
   q             
       �    }          
       
   q      
       
       �    }          
          q      
              �    }                 
   q             
       5�_�   J   L           K   �       ����                                                                                                                                                                                                                                                                                                                                                             f�v     �   �   �   �      ,                            serial_o <= '0';5��    �                    �                    �    �                      �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                 
   �             
       �    �          
          �      
              �    �                 
   �             
       5�_�   K   M           L   �   +    ����                                                                                                                                                                                                                                                                                                                                                             f�     �   �   �   �      .                            parity_bit <= '0';5��    �   +                 �                    5�_�   L   O           M   �   (    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �          )                            word <= data;5��    �                      E      *               5�_�   M   P   N       O   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      ;                        serial_o <= word(signal_bits_sent);5��    �                    �                    �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�   O   Q           P   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      9                        enable <= word(signal_bits_sent);5��    �                    �                    �    �                     �                     �    �                     �                     �    �                     �                     �    �                 
   �             
       �    �   !                  �                     �    �                      �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                 
   �             
       �    �          
       
   �      
       
       �    �          
          �      
              �    �                 
   �             
       5�_�   P   R           Q   �   &    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      =                        shift_data <= word(signal_bits_sent);5��    �   &                  �                     5�_�   Q   S           R   �   &    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      '                        shift_data <= ;5��    �   &                  �                     5�_�   R   T           S   �   '    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      )                        shift_data <= '';5��    �   '                  �                     5�_�   S   U           T   �   '    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �    5��    �                      �                     5�_�   T   V           U   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �                                  5��    �                                          5�_�   U   W           V   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �                                  ''5��    �                                          �    �                                        �    �                     
                     �    �                     	                     �    �                 
                
       �    �   %                                       �    �   $                                       �    �   #                                       �    �   "                                       �    �   !                                       �    �                                           �    �                                          �    �                     
                     �    �                     	                     �    �                 
                
       �    �          
                
              �    �                                        5�_�   V   X           W   �   +    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      +                            shift_data <= 05��    �   *                                       5�_�   W   Y           X   �   *    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      *                            shift_data <= 5��    �   *                                       5�_�   X   Z           Y   �   +    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      ,                            shift_data <= ''5��    �   +                                       5�_�   Y   [           Z   �   -    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      -                            shift_data <= '0'5��    �   -                                       5�_�   Z   \           [   �   !    ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �    �   �   �   �    5��    �                      �              /       5�_�   [   ]           \   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      .                            shift_data <= '0';5��    �                     �                     5�_�   \   ^           ]   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �          .                            shift_data <= '0';5��    �                            /               5�_�   ]   _           ^   �        ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �    �   �   �   �    5��    �                      h              /       5�_�   ^   `           _   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �                              �   �   �   �    5��    �                      2                     �    �                     J                     �    �                     N                     �    �                     M                     �    �                     L                     �    �                     K                     �    �                 
   J             
       �    �          
          J      
              �    �                 
   J             
       5�_�   _   a           `           ����                                                                                                                                                                                                                                                                                                                                                V   !    f�)     �         �    5��                                               5�_�   `   b           a           ����                                                                                                                                                                                                                                                                                                                                                V   !    f�)     �      4   �    �         �    5��                                              5�_�   a   c           b          ����                                                                                                                                                                                                                                                                                                                                                V   !    f�+     �         �      entity shift_reg8 is5��              
          %      
              5�_�   b   d           c   #       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�1     �   "   $   �      &architecture Behavior of shift_reg8 is5��    "          
          �      
              5�_�   c   e           d          ����                                                                                                                                                                                                                                                                                                                                                V   !    f�6     �         �              data: in bit;5��                        b                    5�_�   d   g           e          ����                                                                                                                                                                                                                                                                                                                                                V   !    f�@     �          �      %        q: out bit_vector(7 downto 0)5��                        |                    5�_�   e   h   f       g   $       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�V     �   #   %   �      =   signal vector: bit_vector(7 downto 0) := (others => '0'); 5��    #          )          �      )              5�_�   g   i           h   $       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�Z     �   #   %   �         signal vector: bit; 5��    #                     �                     5�_�   h   j           i   $       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�\     �   #   %   �         signal vector: bit := ; 5��    #                     �                     5�_�   i   l           j   $       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�\     �   #   %   �         signal vector: bit := ''; 5��    #                     �                     5�_�   j   m   k       l   +       ����                                                                                                                                                                                                                                                                                                                                                V   !    f��     �   *   ,   �      &            vector <= (others => '0');5��    *                     0                     5�_�   l   n           m   +       ����                                                                                                                                                                                                                                                                                                                                                V   !    f��     �   *   ,   �                  vector <= ;5��    *                     0                     5�_�   m   o           n   +       ����                                                                                                                                                                                                                                                                                                                                                V   !    f��     �   *   ,   �                  vector <= '';5��    *                     1                     5�_�   n   p           o   -       ����                                                                                                                                                                                                                                                                                                                                                V   !    f��     �   ,   .   �      0            vector <= data & vector(7 downto 1);5��    ,          $          v      $              �    ,                     w                     �    ,                    v                    �    ,                    v                    �    ,                    v                    5�_�   o   q           p   �       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�F     �   �   �   �          parity_bit�   �   �   �              �   �   �   �    5��    �                      k              	       �    �                      k                     �    �                     k              	       �    �                    p                    �    �   	                  u                     �    �                     t                     �    �                     s                     �    �                     r                     �    �                     q                     �    �                    p                    �    �   	                  u                     �    �                     t                     �    �                     s                     �    �                     r                     �    �                     q                     �    �                 
   p             
       �    �                     y                     �    �                     x                     �    �                     w                     �    �   
                  v                     �    �   	                  u                     �    �                     t                     �    �                     s                     �    �                     r                     �    �                     q                     �    �                 
   p             
       �    �          
          p      
              �    �                    p                    �    �                     {                     �    �                     z                     �    �                     y                     �    �                     x                     �    �                     w                     �    �   
                 v                    �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    �    �                    �                     �    �                     �                     �    �   	                 �                    5�_�   p   r           q   �       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�k     �   �   �   �              port map5��    �                     �                     5�_�   q   s           r   �       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�l     �   �   �   �              port map()5��    �                     �                     �    �                 
   �             
       �    �          
          �      
              �    �                    �                    �    �   +                 �                    �    �   +                 �                    �    �   +                 �                    5�_�   r   t           s   ~       ����                                                                                                                                                                                                                                                                                                                                                V   !    f��     �   ~   �   �          �   ~   �   �    5��    ~                      3                     �    ~                     7                     5�_�   s   u           t          ����                                                                                                                                                                                                                                                                                                                                                V   !    f��     �   ~   �   �          signal final_parity5��    ~                     J                     �    ~                    O                    5�_�   t   v           u   �   9    ����                                                                                                                                                                                                                                                                                                                                                V   !    f��     �   �   �   �      :        port map(reset, clock, shift_data, current_parity)5��    �   9                  �                     �    �   ;                 �                    �    �   ;                 �                    �    �   ;                 �                    5�_�   u   w           v   �   H    ����                                                                                                                                                                                                                                                                                                                                                V   !    f��     �   �   �   �      H        port map(reset, clock, shift_data, current_parity, final_parity)5��    �   H                  �                     5�_�   v   x           w   �   -    ����                                                                                                                                                                                                                                                                                                                                                V   !    f��     �   �   �   �                                  �   �   �   �    5��    �                      J                     �    �                     f                     �    �                      j                     �    �                     i                     �    �                     h                     �    �                     g                     �    �                    f                    �    �                    f                    �    �                    f                    �    �   1                  {                     �    �   0                  z                     �    �   /                  y                     �    �   .                 x                    �    �   5                                       �    �   4                  ~                     �    �   3                  }                     �    �   2                  |                     �    �   1                  {                     �    �   0                  z                     �    �   /                  y                     �    �   .              	   x             	       �    �   6                  �                     �    �   5                                       �    �   4                  ~                     �    �   3                  }                     �    �   2                  |                     �    �   1                  {                     �    �   0                  z                     �    �   /                  y                     �    �   .              	   x             	       �    �   .       	          x      	              �    �   .              
   x             
       5�_�   w   y           x   �   .    ����                                                                                                                                                                                                                                                                                                                                                V   !    f�     �   �   �   �      8                            current_parity <= serial_in;5��    �   .       	          x      	              �    �   1                  {                     �    �   0                  z                     �    �   /                  y                     �    �   .              	   x             	       �    �   6                  �                     �    �   5                                       �    �   4                  ~                     �    �   3                  }                     �    �   2                  |                     �    �   1                  {                     �    �   0                  z                     �    �   /                  y                     �    �   .                 x                    �    �   5                                       �    �   4                  ~                     �    �   3                  }                     �    �   2                  |                     �    �   1                  {                     �    �   0                  z                     �    �   /                  y                     �    �   .                 x                    �    �   .                 x                    �    �   .                 x                    �    �   .                 x                    5�_�   x   z           y   �       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�     �   �   �   �      :                            current_parity <= serial_data;5��    �                    f                    �    �                      j                     �    �                     i                     �    �                     h                     �    �                     g                     �    �                    f                    �    �                    f                    �    �                    f                    5�_�   y   {           z   �       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�0     �   �   �   �      8                            final_parity <= serial_data;5��    �                    f                    �    �                     i                     �    �                     h                     �    �                     g                     �    �                    f                    �    �                    f                    �    �                    f                    5�_�   z   |           {   �   )    ����                                                                                                                                                                                                                                                                                                                                                V   !    f�?     �   �   �          :                            current_parity <= serial_data;5��    �                      J      ;               5�_�   {   }           |   �        ����                                                                                                                                                                                                                                                                                                                                                V   !    f�@     �   �   �   �    �   �   �   �    5��    �                      �              ;       5�_�   |   ~           }   �       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�B     �   �   �   �      :                            current_parity <= serial_data;5��    �                     �                     5�_�   }              ~   �   !    ����                                                                                                                                                                                                                                                                                                                                                V   !    f�M     �   �   �          "                        parity_bit5��    �                      m      #               5�_�   ~   �              �   !    ����                                                                                                                                                                                                                                                                                                                                                V   !    f�i     �   �   �   �                                  �   �   �   �    5��    �                      �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    �    �   0                  �                     �    �   /                  �                     �    �   .                 �                    �    �   .                 �                    �    �   .                 �                    �    �   A                  �                     �    �   @                  �                     �    �   ?                 �                    �    �   ?                 �                    �    �   ?                 �                    5�_�      �           �   �   -    ����                                                                                                                                                                                                                                                                                                                                                V   !    f��     �   �   �   �                                  �   �   �   �    5��    �                      g                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                 
   �             
       �    �          
          �      
              �    �                    �                    �    �   ,                  �                     �    �   +                  �                     �    �   *                 �                    �    �   *                 �                    �    �   *                 �                    5�_�   �   �   �       �   �   ?    ����                                                                                                                                                                                                                                                                                                                                                V   !    f��     �   �   �   �      N                            current_parity <= final_parity xor current_parity;5��    �   ?                 �                    �    �   A                  �                     �    �   @                  �                     �    �   ?                 �                    �    �   ?                 �                    �    �   ?                 �                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                V   !    f��    �   �   �          ?                            serial_o <= word(signal_bits_sent);5��    �                      ]      @               5�_�   �   �           �   m       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�     �   n   x   �          �   o   p   �    �   m   p   �          �   m   o   �    5��    m                      !	                     �    m                      !	                     �    m                      !	                     �    m                     !	                     �    n                     &	                    5�_�   �   �           �   o       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�      �   n   p   �      Q        function data_to_parity(data: bit_vector(WIDTH-1 downto 0)) return bit is5��    n                     &	                     5�_�   �   �           �   w        ����                                                                                                                                                                                                                                                                                                                                                V   !    f�(     �   v   w           5��    v                      5
                     5�_�   �   �   �       �   �        ����                                                                                                                                                                                                                                                                                                                                                V   !    f�F     �   �   �              signal final_parity: bit;5��    �                      G                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                                                V   !    f�F     �   �   �              signal current_parity: bit;5��    �                      '                      5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                                                V   !    f�K     �   �   �              parity_process: reg1   I        port map(reset, clock, shift_data, current_parity, final_parity);       5��    �                      `      h               5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V   !    f�N     �                entity reg1 is   
    port (   !        rst, clk, enable: in bit;           d: in bit;           q: out bit       );   end entity;    5��                                v               5�_�   �   �   �       �           ����                                                                                                                                                                                                                                                                                                                                       +           V        f�S     �                 architecture Behavior of reg1 is      signal vector: bit := '0';        begin              process(rst, clk)   	    begin           if rst = '1' then               vector <= '0';   4        elsif rising_edge(clk) and enable = '1' then               vector <= d;           end if;       end process;           q <= vector;          end architecture Behavior;5��                                B              5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                  V        f�T     �                 5��                                               5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �          "                parity_bit <= '1';5��    �                      Q      #               5�_�   �   �   �       �   �        ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �          .                            parity_bit <= '1';5��    �                      �      /               5�_�   �   �   �       �   �   +    ����                                                                                                                                                                                                                                                                                                                                                  V        f�     �   �   �   �      .                            shift_data <= '0';5��    �   +                 1                    5�_�   �   �           �   �   )    ����                                                                                                                                                                                                                                                                                                                                                  V        f�5     �   �   �          *                        shift_data <= '1';5��    �                      �      +               5�_�   �   �           �   �   +    ����                                                                                                                                                                                                                                                                                                                                                  V        f�;     �   �   �          6                        current_parity <= serial_data;5��    �                      �      7               5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                                                  V        f�H     �   �   �          K                            current_parity <= final_parity xor serial_data;5��    �                      ^      L               5�_�   �   �   �       �   �        ����                                                                                                                                                                                                                                                                                                                                                  V        f�`     �   �   �   �      9                            parity_bit <= current_parity;5��    �                    �                    �    �                     �                     �    �                     �                     �    �                 
   �             
       �    �          
          �      
              �    �                    �                    5�_�   �   �           �   �   *    ����                                                                                                                                                                                                                                                                                                                                                  V        f�d     �   �   �   �      *                            shift_data <= 5��    �   *                                       5�_�   �   �           �   �   +    ����                                                                                                                                                                                                                                                                                                                                                  V        f�d     �   �   �   �      ,                            shift_data <= ''5��    �   +                                       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �   �      O                            serial_o <= not data_to_parity(word); -- parity bit5��    �                    G                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �   �      M                            parity <= not data_to_parity(word); -- parity bit5��    �                    G                    �    �                 
   G             
       �    �          
       
   G      
       
       �    �          
          G      
              �    �                 
   G             
       5�_�   �   �           �   �   -    ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �   �      -                            shift_data <= '0'5��    �   -                                       5�_�   �   �           �   �   ,    ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �   �      <                        if stop_bits_sent < (STOP_BITS) then5��    �   ,                 �                    5�_�   �   �           �   �   2    ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �   �      2                        if stop_bits_sent < 2 then5��    �   2                  �                     �    �   6                 �                    5�_�   �   �           �   q       ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   r   t   �          constant STOP_BITS-1�   q   t   �          �   q   s   �    5��    q                                           �    q                                           �    q                                          �    r                                          �    r                     )                     �    r                     (                     �    r                     '                     �    r                     &                     �    r                    %                    �    r                     /                     �    r                     .                     �    r                     -                     �    r                     ,                     �    r                     +                     �    r                     *                     �    r                     )                     �    r                     (                     �    r                     '                     �    r                     &                     �    r                    %                    �    r                    %                    �    r                    %                    �    r                     /                     �    r                    .                    5�_�   �   �           �   |       ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   {   }   �      0        generic map(2+1) -- Stop bits and parity5��    {                                        �    {                                          �    {                                          �    {                 	                	       �    {          	       	         	       	       �    {          	                	              �    {                 	                	       5�_�   �   �           �   �   ,    ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �   �      T                        if stop_bits_sent < 2 then -- numero de stop bits arbitrario5��    �   ,                                     �    �   .                  !                     �    �   -                                        �    �   ,              	                	       �    �   ,       	                	              �    �   ,              	                	       5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                                                  V        f�     �   �   �   �      /                                tx_done <= '1';5��    �                                         5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �          9                            serial_o <= '1'; -- stop bits5��    �                      f      :               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �          #                            -- Data5��    �                      B      $               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �   �      /                            if tx_go = '1' then5��    �                    ~                    �    �   !                  �                     �    �                                           �    �                    ~                    �    �                    ~                    �    �                    ~                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �   �      2                            if starting = '1' then5��    �                    ~                    5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �   �      /                                tx_done <= '0';5��    �                     �                    5�_�   �   �           �   �   #    ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �          0                                serial_o <= '0';5��    �                      �      1               5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �   �    �   �   �   �    5��    �                      �              �       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �          .                            state <= starting;5��    �                      �      /               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �          (                            done <= '0';5��    �                      �      )               5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �           5��    �                      �                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �          &                            -- Control5��    �                      �      '               5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �          0                            start_signal <= '1';5��    �                      �      1               5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �          .                            shift_data <= '1';5��    �                      �      /               5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        f��     �   �   �   �    �   �   �   �    �   �   �          -                                word <= data;5��    �                      P      .               �    �                      P              /       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �           �   -       V        f��     �   �   �   �      .                            shift_data <= '1';5��    �                     l                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �   �    �   �   �   �    5��    �                      �              �       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �          )                state <= idle; -- repouso5��    �                      �      *               5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �   �      0                                serial_o <= '1';5��    �                     �                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �                          done <= '1';5��    �                      �                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �           5��    �                      �                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �                          -- Control5��    �                      �                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �          $                start_signal <= '0';5��    �                      �      %               5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �          "                start_stop <= '0';5��    �                      �      #               5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f��     �   �   �          "                shift_data <= '0';5��    �                      �      #               5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        f��     �   �   �   �    �   �   �   �    �   �   �          8                                word <= (others => '0');5��    �                      �      9               �    �                      �              #       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �           �   !       V        f��     �   �   �   �      "                shift_data <= '0';5��    �                     �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �           �   !       V        f�    �   �   �   �      &                            -- Control5��    �                                          5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                 V       f�S     �   �   �   �      *                                -- Control5��    �           *       &         *       &       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                 V       f�S     �   �   �   �      &                            -- Control5��    �           &       *         &       *       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                 V       f�Z    �          �    �         �    5��                                           )       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                  V       f��     �         �      end architecture Behavior;5��                         <                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                  V       f��    �         �      end architecture ;5��                         ;                     5�_�   �   �           �   j        ����                                                                                                                                                                                                                                                                                                                            a          j          V   *    f�     �   j   l   �    5��    j                      �	                     �    j                      �	                     5�_�   �   �           �   k        ����                                                                                                                                                                                                                                                                                                                            a          j          V   *    f�     �   k   v   �    �   k   l   �    5��    k               
       �	              7      5�_�   �   �           �   l       ����                                                                                                                                                                                                                                                                                                                            a          j          V   *    f�     �   k   m   �          component counter_generic5��    k                    �	                    �    k                     �	                     �    k                     �	                     �    k                 
   �	             
       �    k          
       
   �	      
       
       �    k          
       
   �	      
       
       �    k          
          �	      
              �    k                 
   �	             
       5�_�   �   �           �   m        ����                                                                                                                                                                                                                                                                                                                            m          t   
       V       f�'     �   l   r   �    �   m   n   �    �   l   m                  generic(               MAX_COUNT: natural   
        );           port (   N            clk, rst, start: in bit;                            -- Clock input               done: out bit;   F            count : out natural       -- 6-bit count output (64 steps)   
        );5��    l                      �	                    �    l                      �	              p       5�_�   �   �           �   m       ����                                                                                                                                                                                                                                                                                                                            m          q                 f�*    �   m   r   �      !        rst, clk, enable: in bit;           data: in bit;   %        q: out bit_vector(7 downto 0)       );�   l   n   �      
    port (5��    l                     �	                     �    m                     
                     �    n                     '
                     �    o                     A
                     �    p                     k
                     5�_�   �   �   �       �   �       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    fÊ     �   �   �          .                            shift_data <= '1';5��    �                            /               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    fÌ     �   �   �   �    �   �   �   �    5��    �                      �              /       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    fÍ    �   �   �   �      .                            shift_data <= '1';5��    �                     �                     5�_�   �   �   �       �   �       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f��     �   �   �          .                            shift_data <= '0';5��    �                      �      /               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f��     �   �   �   �                                  �   �   �   �    5��    �                      Z                     �    �                     v                     �    �   !                  {                     �    �                      z                     �    �                    y                    �    �   $                  ~                     �    �   #                  }                     �    �   "                  |                     �    �   !                  {                     �    �                      z                     �    �                    y                    �    �   *                  �                     �    �   )                  �                     �    �   (                  �                     �    �   '                  �                     �    �   &                  �                     �    �   %                                       �    �   $                  ~                     �    �   #                  }                     �    �   "                  |                     �    �   !                  {                     �    �                      z                     �    �                    y                    �    �   #                  }                     �    �   "                  |                     �    �   !                  {                     �    �                      z                     �    �                    y                    �    �   .                  �                     �    �   -                  �                     �    �   ,                  �                     �    �   +                  �                     �    �   *                  �                     �    �   )                  �                     �    �   (                  �                     �    �   '                  �                     �    �   &                  �                     �    �   %                                       �    �   $                  ~                     �    �   #                  }                     �    �   "                  |                     �    �   !                  {                     �    �                      z                     �    �                    y                    �    �                    y                    �    �                    y                    �    �   2                 �                    �    �   6                  �                     �    �   5                  �                     �    �   4                  �                     �    �   3                  �                     �    �   2                 �                    �    �   8                  �                     �    �   7                  �                     �    �   6                  �                     �    �   5                  �                     �    �   4                  �                     �    �   3                  �                     �    �   2                 �                    �    �   2                 �                    �    �   2                 �                    �    �   :                 �                    �    �   :                 �                    �    �   :                 �                    �    �   >                 �                     �    �                      �                     �    �                       �                      5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f��     �   �   �   �    �   �   �   �    5��    �                      �              /       5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f��     �   �   �           5��    �                      �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f��     �   �   �   �      .                            shift_data <= '0';5��    �                     �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f��    �   �   �   �                                       �   �   �   �    5��    �                      �              !       �    �                      �                     �    �                      �                     �    �                      �                     �    �   "                 �                    5�_�   �   �   �       �   �       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f�{     �   �   �   �                                  �   �   �   �    5��    �                      �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    �    �   .                                       �    �   -                                     �    �   -                                     �    �   -                                     5�_�   �   �           �   �   1    ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    fȃ    �   �   �   �      1                            parallel_data <= word5��    �   1                                       5�_�   �   �           �   H       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f�O    �   G   I   �      entity serial_in is5��    G                                          5�_�   �   �           �   V   $    ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f�f    �   U   W   �      'architecture Behavioral of serial_in is5��    U   $                  �                     5�_�   �   �   �       �   C       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f��     �   C   E   �    5��    C                      �                     5�_�   �   �           �   D        ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f��    �   D   a   �    �   D   E   �    5��    D                      �              7      5�_�   �   �           �   Q       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f�	     �   P   R   �      )    signal counter: unsigned(9 downto 0);5��    P                    �                    5�_�   �   �           �   Q       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f�     �   P   R   �      )    signal counter: unsigned(2 downto 0);5��    P                    �                    5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f�     �   Y   [   �      *            if counter = "1111111111" then5��    Y          
          �      
              5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f�i     �   �   �   �          �   �   �   �    5��    �                      �                     �    �                      �                     �    �                      �                     �    �                     �                     �    �                     �                     �    �   	                  �                     �    �                     �                     �    �                     �                     �    �                     �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f�n     �   �   �              si5��    �                      �                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f�o     �   �   �           5��    �                      �                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �           ~           V        f�{     �   �   �   �    5��    �                                           �    �                                           5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �           ~           V        f�{     �   �   �   �    �   �   �   �    5��    �               
       	              7      5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �           ~           V        f�}     �   �   �   �          component counter_generic5��    �                                        �    �                                          �    �                                          �    �                                          �    �                                        �    �                                        �    �                                        5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �   
       V       fۊ     �   �   �   �    �   �   �   �    �   �   �                  generic(               MAX_COUNT: natural   
        );           port (   N            clk, rst, start: in bit;                            -- Clock input               done: out bit;   F            count : out natural       -- 6-bit count output (64 steps)   
        );5��    �                                           �    �                                     C       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 fێ     �   �   �   �              clk_in: in bit;           clk_out: out bit       );�   �   �   �      
    port (5��    �                     $                     �    �                     3                     �    �                     O                     �    �                     l                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 fۖ     �   �   �   �              port�   �   �   �          clocking: slow_clk�   �   �   �          �   �   �   �    5��    �                      �                     �    �                      �                     �    �                      �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    �    �                    �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 fۭ     �   �   �   �              port map5��    �                     �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 fۮ     �   �   �   �              port map()5��    �                     �                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 f۵     �   �   �   �               port map(clock, new_clk)5��    �                                           5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 f۷     �   �   �   �          �   �   �   �    5��    �                      �                     �    �                     �                     �    �                 
   �             
       �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      F        port map(clock, reset, start_stop, done_stop, stop_bits_sent);5��    �                                        �    �                                          �    �                                          �    �                                          �    �                                        �    �                                        �    �                                        5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      >        port map(reset, clock, shift_data, serial_data, word);5��    �                    �                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      <        port map(reset, new, shift_data, serial_data, word);5��    �                     �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      >        port map(reset, new[], shift_data, serial_data, word);5��    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �   �       �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �      "        if rising_edge(clock) then5��    �                    �                    �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f�     �   �   �   �      $        if rising_edge(new_clk) then5��    �                    �                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f�8    �   �   �   �      "        if rising_edge(clock) then5��    �                    �                    �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   s   $    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�a     �   r   t   �      )architecture Behavioral of serial_in_V is5��    r   $                  �	                     5�_�   �   �           �   s   $    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�a     �   r   t   �      (architecture Behavioral of serial_inV is5��    r   $                  �	                     5�_�   �   �           �   e       ����                                                                                                                                                                                                                                                                                                                            �          �                 f�k     �   d   f   �      entity serial_in_V is5��    d                     O                     5�_�   �   �           �   e       ����                                                                                                                                                                                                                                                                                                                            �          �                 f�l    �   d   f   �      entity serial_inis5��    d                     O                     5�_�   �   �           �   Q   (    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�B     �   P   R   �      )    signal counter: unsigned(1 downto 0);5��    P   (                  �                     5�_�   �              �   Q   ,    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�F     �   P   R   �      -    signal counter: unsigned(1 downto 0) := ;5��    P   ,                  �                     5�_�   �                Q   -    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�G     �   P   R   �      /    signal counter: unsigned(1 downto 0) := '';5��    P   ,                  �                     �    P   ,                  �                     5�_�                  Q   ,    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�G     �   P   R   �      -    signal counter: unsigned(1 downto 0) := ;5��    P   ,                  �                     5�_�                 Q   -    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�H     �   P   R   �      /    signal counter: unsigned(1 downto 0) := "";5��    P   -                  �                     5�_�                 [       ����                                                                                                                                                                                                                                                                                                                            �          �                 f�     �   Z   \   �      -                clk_out <= not current_state;5��    Z                    �                    �    Z                     �                     �    Z                     �                     �    Z                    �                    �    Z                    �                    �    Z                    �                    5�_�                 ^       ����                                                                                                                                                                                                                                                                                                                            �          �                 f�!    �   _   a   �          clk_out�   ^   a   �          �   ^   `   �    5��    ^                                           �    ^                                           �    ^                                          �    _                                          �    _                                          �    _                                          �    _                                          �    _                                        �    _                                        �    _                                        �    _                                          �    _                                          �    _                                          �    _                                        �    _                                        �    _                                        5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f�x    �   �   �   �          process(clock) is5��    �                    �                    �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�                 g       ����                                                                                                                                                                                                                                                                                                                            �          �                 f�B    �   f   h   �      entity serial_in is5��    f                     |                     �    f                    |                    5�_�                 u   $    ����                                                                                                                                                                                                                                                                                                                            �          �                 f��    �   t   v   �      'architecture Behavioral of serial_in is5��    t   $                  �	                     5�_�    	             g       ����                                                                                                                                                                                                                                                                                                                            �          �                 f�u     �   f   h   �      entity serial_inV is5��    f                     |                     5�_�    
          	   u   $    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�y    �   t   v   �      (architecture Behavioral of serial_inv is5��    t   $                  �	                     5�_�  	            
   Z       ����                                                                                                                                                                                                                                                                                                                            �          �                 f�     �   Y   [   �      "            if counter = "11" then5��    Y                    �                    5�_�  
               Q       ����                                                                                                                                                                                                                                                                                                                            �          �                 f�     �   P   R   �      1    signal counter: unsigned(1 downto 0) := "00";5��    P                    �                    5�_�                 Q   -    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�    �   P   R   �      1    signal counter: unsigned(0 downto 0) := "00";5��    P   -                  �                     5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��    �   �   �   �      L        port map(clock, reset, start_signal, done_signal, signal_bits_sent);5��    �                    �                    �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �          *                        shift_data <= '1';5��    �                      �      +               5�_�                 �        ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �    �   �   �   �    5��    �                      <              +       5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��    �   �   �   �      *                        shift_data <= '1';5��    �                     T                     5�_�               �   1    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�     �   �   �                                     �   �   �   �    5��    �                      N                     �    �                     j                     �    �                     l                     �    �                     k                     �    �                    j                    �    �                    j                    �    �                 	   j             	       �    �   $                  r                     5�_�                 �   $    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�     �   �   �         $                            done <= 5��    �   $                  r                     5�_�                 �   %    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�     �   �   �         &                            done <= ''5��    �   %                  s                     5�_�                 �   '    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�     �   �   �         '                            done <= '1'5��    �   '                  u                     5�_�                 �        ����                                                                                                                                                                                                                                                                                                                            �   '       �   #       V   '    f��    �   �   �          B                            if stop_bits_sent = (STOP_BITS-1) then   ,                                done <= '1';   #                            end if;5��    �                      x      �               5�_�               �   *    ����                                                                                                                                                                                                                                                                                                                            �   '       �   #       V   '    f��     �   �   �   �      /                            if start = '1' then5��    �   *                  �                     �    �   -                  �                     �    �   ,                  �                     �    �   +                 �                    �    �   5                  �                     �    �   4                  �                     �    �   3                  �                     �    �   2                  �                     �    �   1                  �                     �    �   0                  �                     �    �   /                  �                     �    �   .                  �                     �    �   -                  �                     �    �   ,                  �                     �    �   +                 �                    �    �   +                 �                    �    �   +                 �                    5�_�                 �   9    ����                                                                                                                                                                                                                                                                                                                            �   '       �   #       V   '    f��     �   �   �   �      >                            if start = '1' serial_data =  then5��    �   9                  �                     5�_�                 �   :    ����                                                                                                                                                                                                                                                                                                                            �   '       �   #       V   '    f��     �   �   �   �      @                            if start = '1' serial_data = '' then5��    �   :                  �                     5�_�                 �   *    ����                                                                                                                                                                                                                                                                                                                            �   '       �   #       V   '    f��     �   �   �   �      A                            if start = '1' serial_data = '0' then5��    �   *                  �                     5�_�                 �   &    ����                                                                                                                                                                                                                                                                                                                            �   '       �   #       V   '    f�     �   �   �   �      +                        if start = '1' then5��    �   &                  �                     �    �   -                  �                     �    �   ,                  �                     �    �   +                 �                    �    �   +                 �                    �    �   +                 �                    5�_�                  �   9    ����                                                                                                                                                                                                                                                                                                                            �   '       �   #       V   '    f�     �   �   �   �      >                        if start = '1' and serial_data =  then5��    �   9                  �                     5�_�                    �   :    ����                                                                                                                                                                                                                                                                                                                            �   '       �   #       V   '    f�     �   �   �   �      @                        if start = '1' and serial_data = '' then5��    �   :                  �                     5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �   '       �   #       V   '    f�     �   �   �   �                      done <= '0';5��    �                    �                    5�_�               g       ����                                                                                                                                                                                                                                                                                                                            �          �                 f�     �   f   h   �      entity serial_inv is5��    f                     z                     5�_�                 u   $    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�    �   t   v   �      (architecture Behavioral of serial_inv is5��    t   $                  �	                     5�_�                   u   $    ����                                                                                                                                                                                                                                                                                                                            �          �                 f�     �   t   v   �      'architecture Behavioral of serial_in is5��    t   $                  �	                     5�_�   �           �   �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f��     �   �   �   �          process() is5��    �                     �                     5�_�   �           �   �   C       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f��     �   C   D   �    �   C   D   �      library IEEE;   use IEEE.NUMERIC_BIT.all;       entity slow_clk is   
    port (           clk_in: in bit;           clk_out: out bit       );   end entity slow_clk;       architecture rtl of slow_clk is       )    signal counter: unsigned(9 downto 0);   (    signal current_state: bit := clk_in;          begin              timing: process(clk_in)   	    begin   #        if rising_edge(clk_in) then   #            counter <= counter + 1;   *            if counter = "1111111111" then   -                clk_out <= not current_state;               end if;           end if;       end process timing;          end architecture rtl;5��    C                      �              7      5�_�   �           �   �   �       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f�k     �   �   �   �      T                            parallel_data <= not data_to_parity(word); -- parity bit5��    �          
          �      
              �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �           �   �   �       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f�!     �   �   �        5��    �                            v               5�_�   �   �   �   �   �   �        ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f     �   �   �   �    �   �   �   �      B                            if stop_bits_sent = (STOP_BITS-1) then   ,                                done <= '1';   #                            end if;5��    �                      ^              �       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f     �   �   �   �      D                            if signal_bits_sent = (STOP_BITS-1) then5��    �                    }                    �    �   "                  �                     �    �   !                                       �    �                      ~                     �    �                    }                    �    �                    }                    �    �                    }                    �    �                    }                    5�_�   �   �           �   �   3    ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f     �   �   �   �      @                            if signal_bits_sent = (WIDTH-1) then5��    �   3       	          �      	              �    �   4                  �                     �    �   3                 �                    �    �   3                 �                    �    �   3                 �                    �    �   3                 �                    5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f     �   �   �   �      2                                shift_data <= '1';5��    �                     �                    �    �   "                  �                     �    �   !                  �                     �    �                  
   �             
       �    �   )                  �                     �    �   (                  �                     �    �   '                  �                     �    �   &                  �                     �    �   %                  �                     �    �   $                  �                     �    �   #                  �                     �    �   "                  �                     �    �   !                  �                     �    �                  
   �             
       �    �           
       
   �      
       
       �    �           
          �      
              �    �                  
   �             
       5�_�   �   �           �   �   /    ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f   	 �   �   �   �      2                                shift_data <= '0';5��    �   /                 �                    5�_�   �               �   �   -    ����                                                                                                                                                                                                                                                                                                                            �   +       �   #       V   +    f¶   
 �   �   �        5��    �                      q      /               5�_�   �           �   �   �   +    ����                                                                                                                                                                                                                                                                                                                            m          q                 f�p     �   �   �   �       5��    �                      �              !       �    �                       �                      5�_�   �           �   �   �        ����                                                                                                                                                                                                                                                                                                                                                  V        f�_     �   �   �        5��    �                      �      :               5�_�   �           �   �   �        ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �        5��    �                            /               5�_�   �           �   �   �        ����                                                                                                                                                                                                                                                                                                                                                  V        f��     �   �   �        5��    �                      �      /               5�_�   �           �   �           ����                                                                                                                                                                                                                                                                                                                                                V   !    f�O     �              5��                                A               5�_�   �           �   �   �        ����                                                                                                                                                                                                                                                                                                                                                V   !    f�>     �   �   �        5��    �                      �      h               5�_�   �           �   �   �   5    ����                                                                                                                                                                                                                                                                                                                                                V   !    f��     �   �   �   �      ;                        current_parity <= serial_data xor ;5��    �   5                  �                     5�_�   j           l   k   $       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�f     �   #   %   �         signal vector: bit; 5��    #                     �                     5�_�   e           g   f   $       ����                                                                                                                                                                                                                                                                                                                                                V   !    f�O     �   #   %        5��    #                      �      >               5�_�   M           O   N   �       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   �   �   �      9                        enable <= word(signal_bits_sent);5��    �                    �                    �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�                             ����                                                                                                                                                                                                                                                                                                                                                             fM^     �         �       �         �           �         �    �         �      !e n t i t y s e r i a l _ i n i s   g en e r ic (   POLARITY : boolean := TRUE;   WIDTH: n a t u r a l := 8 ;   PARITY : n a t u r a l := 1 ;   CLOCK_MUL: p o s i t i v e := 4   ) ;   po r t (   Bclock , r e s e t , s t a r t , s e r i a l _ d a t a : in b i t ;   (done , p a r i t y _ b i t : out b i t ;   Hp a r a l l e l _ d a t a : out b i t _ v e c t o r (WIDTH−1 downto 0)   ) ;   end s e r i a l _ i n ;5��                          >                     �                          >                     �                         ?              �      5��