Vim�UnDo� �w^�qKw�މX{��U����c���a�   �        �                          f(l�    _�                             ����                                                                                                                                                                                                                                                                                                                                                  V        f(J     �                 library IEEE;   use IEEE.NUMERIC_BIT.all;       entity reg32 is   
    port (   !        rst, clk, enable: in bit;   )        init: in bit_vector(31 downto 0);   &        d: in bit_vector(31 downto 0);   &        q: out bit_vector(31 downto 0)       );   end entity reg32;       !architecture Behavior of reg32 is   *    signal value: bit_vector(31 downto 0);   begin              process(rst, clk)   	    begin           if rst = '1' then               value <= init;   4        elsif rising_edge(clk) and enable = '1' then               value <= D;           end if;       end process;           q <= value;          end architecture Behavior;    5��                                   E              5�_�                            ����                                                                                                                                                                                                                                                                                                                                       !           V        f(J#     �              !   library IEEE;   use IEEE.NUMERIC_BIT.all;       entity shift_reg512 is   
    port (   !        rst, clk, enable: in bit;   )        data: in bit_vector(31 downto 0);   '        d: in bit_vector(511 downto 0);   '        q: out bit_vector(511 downto 0)       );   end entity shift_reg512;       (architecture Behavior of shift_reg512 is   ,   signal vector: bit_vector(511 downto 0);        begin              process(rst, clk)   	    begin           if rst = '1' then               vector <= d;   4        elsif rising_edge(clk) and enable = '1' then   2            vector <= vector(479 downto 0) & data;           end if;       end process;           q <= vector;          end architecture Behavior;       library IEEE;   use IEEE.NUMERIC_BIT.ALL;    5��            !                       �              5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �                   V       f(J)     �   �   �          entity adder32 is   port(   &    a, b : in bit_vector(31 downto 0);   #    s : out bit_vector(31 downto 0)       );   end adder32;       %architecture behavioral of adder32 is   +    signal carry : bit_vector(31 downto 0);   begin   "    sum: for i in 0 to 30 generate   +        s(i) <= A(i) xor B(i) xor carry(i);   T        carry(i+1) <= (A(i) and B(i)) or (A(i) and carry(i)) or (B(i) and carry(i));       end generate;       +    s(31) <= A(31) xor B(31) xor carry(31);         end behavioral;5��    �                             �              5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f(J*    �   �   �           5��    �                                           5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f(J4    �   �   �              -- process(clk, rst)       -- begin       --     if rst = '1' then       --         enable <= '1';   &    --     elsif rising_edge(clk) then   %    --         if iteration = 63 then   !    --             enable <= '0';       --         end if;       --       --     end if;       --       -- end process;    5��    �                      �                    5�_�                            ����                                                                                                                                                                                                                                                                                                                                       �           V        f(l�     �       #          entity multisteps is�              �             �   
    port (   !        clk, rst, enable: in bit;   +        msgi : in bit_vector(511 downto 0);   ,        haso : out bit_vector(255 downto 0);           done : out bit       );   end multisteps;       !architecture rtl of multisteps is           component stepfun  is           port (   D        	ai, bi, ci, di, ei, fi, gi, hi: in bit_vector(31 downto 0);   ,            kpw: in bit_vector(31 downto 0);   G            ao, bo, co, do, eo, fo, go, ho: out bit_vector(31 downto 0)   
        );       end component;           component reg32 is           port (   %            rst, clk, enable: in bit;   -            init: in bit_vector(31 downto 0);   *            d: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           component shift_reg512 is           port (   %            rst, clk, enable: in bit;   -            data: in bit_vector(31 downto 0);   +            d: in bit_vector(511 downto 0);   +            q: out bit_vector(511 downto 0)   
        );       end component;       !    component counter_generic  is           generic(               MAX_COUNT: natural   
        );           port (   N            clk, rst, start: in bit;                            -- Clock input               done: out bit;   F            count : out natural       -- 6-bit count output (64 steps)   
        );       end component;           component adder32  is           port (   +            a : in bit_vector(31 downto 0);   +            b : in bit_vector(31 downto 0);   +            s : out bit_vector(31 downto 0)   
        );       end component;           component sigma0 is            port(   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;              component sigma1 is           port(   *            x: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           -- Constants   9    constant h0 : bit_vector(31 downto 0) := x"6a09e667";   9    constant h1 : bit_vector(31 downto 0) := x"bb67ae85";   9    constant h2 : bit_vector(31 downto 0) := x"3c6ef372";   9    constant h3 : bit_vector(31 downto 0) := x"a54ff53a";   9    constant h4 : bit_vector(31 downto 0) := x"510e527f";   9    constant h5 : bit_vector(31 downto 0) := x"9b05688c";   9    constant h6 : bit_vector(31 downto 0) := x"1f83d9ab";   9    constant h7 : bit_vector(31 downto 0) := x"5be0cd19";           -- Signals   C    type aux_signals is array (0 to 63) of bit_vector(31 downto 0);        signal k_const: aux_signals;           signal iteration: natural;       signal ended: bit;   +    signal w_vec: bit_vector(511 downto 0);   +    signal next_w: bit_vector(31 downto 0);   .    signal current_w: bit_vector(31 downto 0);   .    signal current_k: bit_vector(31 downto 0);   0    signal current_kpw: bit_vector(31 downto 0);       7    signal op1, op2, op3, op4: bit_vector(31 downto 0);   '    signal av: bit_vector(31 downto 0);   '    signal bv: bit_vector(31 downto 0);   '    signal cv: bit_vector(31 downto 0);   '    signal dv: bit_vector(31 downto 0);   '    signal ev: bit_vector(31 downto 0);   '    signal fv: bit_vector(31 downto 0);   '    signal gv: bit_vector(31 downto 0);   '    signal hv: bit_vector(31 downto 0);   *    signal a_reg: bit_vector(31 downto 0);   *    signal b_reg: bit_vector(31 downto 0);   *    signal c_reg: bit_vector(31 downto 0);   *    signal d_reg: bit_vector(31 downto 0);   *    signal e_reg: bit_vector(31 downto 0);   *    signal f_reg: bit_vector(31 downto 0);   *    signal g_reg: bit_vector(31 downto 0);   *    signal h_reg: bit_vector(31 downto 0);       begin              -- Assynchronous operations       k_const(0) <= x"428a2f98";       k_const(1) <= x"71374491";       k_const(2) <= x"b5c0fbcf";       k_const(3) <= x"e9b5dba5";       k_const(4) <= x"3956c25b";       k_const(5) <= x"59f111f1";       k_const(6) <= x"923f82a4";       k_const(7) <= x"ab1c5ed5";       k_const(8) <= x"d807aa98";       k_const(9) <= x"12835b01";       k_const(10) <= x"243185be";       k_const(11) <= x"550c7dc3";       k_const(12) <= x"72be5d74";       k_const(13) <= x"80deb1fe";       k_const(14) <= x"9bdc06a7";       k_const(15) <= x"c19bf174";       k_const(16) <= x"e49b69c1";       k_const(17) <= x"efbe4786";       k_const(18) <= x"0fc19dc6";       k_const(19) <= x"240ca1cc";       k_const(20) <= x"2de92c6f";       k_const(21) <= x"4a7484aa";       k_const(22) <= x"5cb0a9dc";       k_const(23) <= x"76f988da";       k_const(24) <= x"983e5152";       k_const(25) <= x"a831c66d";       k_const(26) <= x"b00327c8";       k_const(27) <= x"bf597fc7";       k_const(28) <= x"c6e00bf3";       k_const(29) <= x"d5a79147";       k_const(30) <= x"06ca6351";       k_const(31) <= x"14292967";       k_const(32) <= x"27b70a85";       k_const(33) <= x"2e1b2138";       k_const(34) <= x"4d2c6dfc";       k_const(35) <= x"53380d13";       k_const(36) <= x"650a7354";       k_const(37) <= x"766a0abb";       k_const(38) <= x"81c2c92e";       k_const(39) <= x"92722c85";       k_const(40) <= x"a2bfe8a1";       k_const(41) <= x"a81a664b";       k_const(42) <= x"c24b8b70";       k_const(43) <= x"c76c51a3";       k_const(44) <= x"d192e819";       k_const(45) <= x"d6990624";       k_const(46) <= x"f40e3585";       k_const(47) <= x"106aa070";       k_const(48) <= x"19a4c116";       k_const(49) <= x"1e376c08";       k_const(50) <= x"2748774c";       k_const(51) <= x"34b0bcb5";       k_const(52) <= x"391c0cb3";       k_const(53) <= x"4ed8aa4a";       k_const(54) <= x"5b9cca4f";       k_const(55) <= x"682e6ff3";       k_const(56) <= x"748f82ee";       k_const(57) <= x"78a5636f";       k_const(58) <= x"84c87814";       k_const(59) <= x"8cc70208";       k_const(60) <= x"90befffa";       k_const(61) <= x"a4506ceb";       k_const(62) <= x"bef9a3f7";       k_const(63) <= x"c67178f2";           -- W combinational   <    int1: sigma1 port map(w_vec(63 downto 32), op1); -- t-14   =    int2: sigma0 port map(w_vec(479 downto 448), op2); -- t-1   *    int4: adder32 port map(op1, op2, op3);   [    int3: adder32 port map(w_vec(223 downto 192), w_vec(511 downto 480), op4); -- t-9 and t   -    int5: adder32 port map(op3, op4, next_w);           -- W sequential   L    shf_w: shift_reg512 port map (rst, clk, not ended, next_w, msgi, w_vec);       B    get_kpw: adder32 port map (current_w, current_k, current_kpw);           counter: counter_generic            generic map(64)   6        port map (clk, rst, enable, ended, iteration);       D    a_register: reg32 port map (rst, clk, not ended, h0, av, a_reg);   D    b_register: reg32 port map (rst, clk, not ended, h1, bv, b_reg);   D    c_register: reg32 port map (rst, clk, not ended, h2, cv, c_reg);   D    d_register: reg32 port map (rst, clk, not ended, h3, dv, d_reg);   D    e_register: reg32 port map (rst, clk, not ended, h4, ev, e_reg);   D    f_register: reg32 port map (rst, clk, not ended, h5, fv, f_reg);   D    g_register: reg32 port map (rst, clk, not ended, h6, gv, g_reg);   D    h_register: reg32 port map (rst, clk, not ended, h7, hv, h_reg);       >    get_aout: adder32 port map (h0, a_reg, haso(31 downto 0));   ?    get_bout: adder32 port map (h1, b_reg, haso(63 downto 32));   ?    get_cout: adder32 port map (h2, c_reg, haso(95 downto 64));   @    get_dout: adder32 port map (h3, d_reg, haso(127 downto 96));   A    get_eout: adder32 port map (h4, e_reg, haso(159 downto 128));   A    get_fout: adder32 port map (h5, f_reg, haso(191 downto 160));   A    get_gout: adder32 port map (h6, g_reg, haso(223 downto 192));   A    get_hout: adder32 port map (hv, h_reg, haso(255 downto 224));           step: stepfun port map (           ai => a_reg,           bi => b_reg,           ci => c_reg,           di => d_reg,           ei => e_reg,           fi => f_reg,           gi => g_reg,           hi => h_reg,           kpw => current_kpw,           ao => av,           bo => bv,           co => cv,           do => dv,           eo => ev,           fo => fv,           go => gv,           ho => hv       );           done <= ended;   '    current_w <= w_vec(511 downto 480);   $    current_k <= k_const(iteration);          end architecture rtl;5��           �                      �              �                                                  �                    !                             5�_�                             ����                                                                                                                                                                                                                                                                                                                                       "           V        f(l�    �   �                �   �            �                  library IEEE;�               �             !   use IEEE.NUMERIC_BIT.ALL;       entity counter_6bit is   
    port (   C        clk, rst: in bit;                            -- Clock input           done: out bit;   O        count : out unsigned(5 downto 0)       -- 6-bit count output (64 steps)       );   end counter_6bit;       #architecture rtl of counter_6bit is   )    signal counter: unsigned(5 downto 0);       begin              counting: process(clk, rst)   	    begin           if rst = '1' then   '            counter <= (others => '0');               done <= '0';   #        elsif rising_edge(clk) then   ,            if to_integer(counter) = 63 then                   done <= '1';               else   '                counter <= counter + 1;               end if;           end if;       end process counting;           count <= counter;          end architecture rtl;    5��           !                      �              �                                                  �                    �                      �      �    �              f       �              �      5��