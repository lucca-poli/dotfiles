Vim�UnDo� h���� 룡�����A�b��EWX����A�   D   n	constant asserts: DwordArray(test_size - 1 downto 0) := (x"DA5698BE", x"DA5698BE", x"B8A4E897", x"27D75F9C");   "   F                           fm   	 _�                         !    ����                                                                                                                                                                                                                                                                                                                                                             f�    �      !   ?      #	constant test_size: positive := 4;5��       !                                     5�_�                   7   
    ����                                                                                                                                                                                                                                                                                                                            7          7   
       v       f��    �   6   8   ?      			assert check = asserts(i)5��    6   
                 �                    5�_�                   7   
    ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f�_     �   6   8   ?      			assert false5��    6   
                 �                    5�_�      	              7       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f�e     �   6   8   ?      			assert check = asserts5��    6                     �                     5�_�      
           	   7       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f�e     �   6   8   ?      			assert check = asserts()5��    6                     �                     5�_�   	              
   9       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f�y     �   9   ;   ?    �   9   :   ?    5��    9                      q              �       5�_�   
                 :       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f��     �   9   ;   @      �				report "Entrada: " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    9                    }                    �    9                    �                    5�_�                    :       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f��     �   9   ;   @      �				report "haso0 : " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    9                     �                     5�_�                    :   ,    ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f��     �   9   ;   @      �				report "haso0: " &  to_hstring(unsigned(datas(i))) & " Esperado: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    9   ,                 �                    5�_�                    :   8    ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f��     �   9   ;   @      �				report "haso0: " &  to_hstring(unsigned(check)) & " Esperado: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    9   8                 �                    5�_�                    :   ^    ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f��     �   9   ;   @      �				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada: " & to_hstring(unsigned(asserts(i))) & " Recebido: " & to_hstring(unsigned(check))5��    9   ^                 �                    5�_�                    :   h    ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f��     �   9   ;   @      �				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada: " & to_hstring(unsigned(datas(i))) & " Recebido: " & to_hstring(unsigned(check))5��    9   h       .           �      .               5�_�                    :   h    ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f��     �   9   ;   @      h				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada: " & to_hstring(unsigned(datas(i)))5��    9   h                  �                     5�_�                    ;       ����                                                                                                                                                                                                                                                                                                                            :   h       7          V   t    f��    �   ;   @   @    �   ;   <   @    5��    ;                      �              4      5�_�                    ?   D    ����                                                                                                                                                                                                                                                                                                                            :   h       7          V   t    f��    �   >   @   D      i				report "haso0: " &  to_hstring(unsigned(check)) & " para entrada: " & to_hstring(unsigned(datas(i)));5��    >   D                                       5�_�                    4       ����                                                                                                                                                                                                                                                                                                                                                             f
�     �   3   5   D      			wait for 4*half_period;5��    3                    h                    5�_�                    ;       ����                                                                                                                                                                                                                                                                                                                                                             f
�    �   :   <   D      			wait for 4*half_period;5��    :                    �                    5�_�                    !   =    ����                                                                                                                                                                                                                                                                                                                            !   7       !   <       v   ?    fK     �       "   D      L	constant datas: ByteArray(test_size - 1 downto 0) := (x"00", x"01", x"02");5��        =                  Q                     5�_�                    !   =    ����                                                                                                                                                                                                                                                                                                                            !   7       !   <       v   ?    fK     �       "   D      M	constant datas: ByteArray(test_size - 1 downto 0) := (x"00",  x"01", x"02");�   !   "   D    5��        >                  R                     5�_�                   "   F    ����                                                                                                                                                                                                                                                                                                                            "   F       "   :       v   =    fU    �   !   #   D      a	constant asserts: DwordArray(test_size - 1 downto 0) := (x"DA5698BE", x"B8A4E897", x"27D75F9C");�   "   #   D    5��    !   G                  �                     5�_�                        "    ����                                                                                                                                                                                                                                                                                                                            "   F       "   :       v   =    fd    �      !   D      #	constant test_size: positive := 3;5��       !                                     5�_�                   !   >    ����                                                                                                                                                                                                                                                                                                                            !   >       !   D       v   G    fV     �       "   D      S	constant datas: ByteArray(test_size - 1 downto 0) := (x"00", x"00", x"01", x"02");5��        >                  R                     5�_�                   !   D    ����                                                                                                                                                                                                                                                                                                                            !   >       !   D       v   G    fY     �       "   D      L	constant datas: ByteArray(test_size - 1 downto 0) := (x"00", x"01", x"02");�   !   "   D    5��        E                  Y                     5�_�                     "   F    ����                                                                                                                                                                                                                                                                                                                            "   F       "   R       v   U    fj     �   !   #   D      n	constant asserts: DwordArray(test_size - 1 downto 0) := (x"DA5698BE", x"DA5698BE", x"B8A4E897", x"27D75F9C");5��    !   F                  �                     5�_�                      "   R    ����                                                                                                                                                                                                                                                                                                                            "   F       "   R       v   U    fl   	 �   !   #   D      a	constant asserts: DwordArray(test_size - 1 downto 0) := (x"DA5698BE", x"B8A4E897", x"27D75F9C");�   "   #   D    5��    !   S                  �                     5�_�                    !   C    ����                                                                                                                                                                                                                                                                                                                            !   >       !   D       v   G    fW     �   !   "   D    �       "   D      S	constant datas: ByteArray(test_size - 1 downto 0) := (x"00", x"01",x"00",  x"02");5��        D                  X                     5�_�                    !   >    ����                                                                                                                                                                                                                                                                                                                            !   >       !   C       v   F    fP     �       "   D      M	constant datas: ByteArray(test_size - 1 downto 0) := (x"00",  x"01", x"02");5��        >                  R                     5�_�                    "   E    ����                                                                                                                                                                                                                                                                                                                            "   F       "   :       v   =    fS     �   "   #   D    �   !   #   D      n	constant asserts: DwordArray(test_size - 1 downto 0) := (x"DA5698BE",x"DA5698BE",  x"B8A4E897", x"27D75F9C");5��    !   F                  �                     5�_�                   4       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f�$     �   3   5   ?      			wait until rising_edge;5��    3                    d                    �    3                    h                    �    3                     l                     �    3                     k                     �    3                    j                    �    3                    j                    �    3                    j                    5�_�                    4       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f�)     �   3   5   ?      			wait until rising_edge();5��    3                     u                     5�_�                     4       ����                                                                                                                                                                                                                                                                                                                            4          4          v   !    f�)     �   3   5   ?       			wait until rising_edge(done);5��    3                     v                     5�_�                    8       ����                                                                                                                                                                                                                                                                                                                                                V   &    f�Z     �   8   9   ?    �   8   9   ?      use std.textio.all;5��    8                      ^                     5��