Vim�UnDo� �L LT��O��㠍o��H}��!Oo�   g   !architecture rtl of serial_out is   4                      f�    _�                        #    ����                                                                                                                                                                                                                                                                                                                                                             f�    �         o      /        data : in bit_vector(WIDTH-1 downto 0);5��       "                 o                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f�     �         o    �         o    5��                                               5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             f�     �                 -- Transmissao serial:5��                                                  5�_�                       
    ����                                                                                                                                                                                                                                                                                                                                                             f�     �          �      entity reg32 is5��        
                 
                     5�_�                            ����                                                                                                                                                                                                                                                                                                                               
                 V   
    f�     �   
             *    signal value: bit_vector(31 downto 0);�                &        q: out bit_vector(31 downto 0)�                &        d: in bit_vector(31 downto 0);�         �      )        init: in bit_vector(31 downto 0);5��                        X                     �                        ~                     �                        �                     �    
                    
                    5�_�                           ����                                                                                                                                                                                                                                                                                                                               
                 V   
    f�     �      	   �      end entity reg32;5��                        �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                               
                 V   
    f�     �          �      entity reg8 is5��        
                  
                      5�_�      	                 
    ����                                                                                                                                                                                                                                                                                                                               
                 V   
    f�     �          �      entity reg is5��                                              �                                              �                                              �                                              5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                               
                 V   
    f�     �      	   �      end entity reg8;5��                        �                     �                         �                      �                        �                     �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     �                        �                     �                        �                     �                        �                     5�_�   	              
   
       ����                                                                                                                                                                                                                                                                                                                               
                 V   
    f�     �   	      �      !architecture Behavior of reg32 is5��    	                    �                     �    	                    �                     �    	                    �                     �    	                    �                     5�_�   
                         ����                                                                                                                                                                                                                                                                                                                                       &          V   #    f
     �      	   �    �         �    5��                                         �       5�_�                           ����                                                                                                                                                                                                                                                                                                                            '          -          V   #    f     �                #        POLARITY : boolean := TRUE;5��                          #       $               5�_�                           ����                                                                                                                                                                                                                                                                                                                            &          ,          V   #    f     �                        PARITY : natural := 1 ;5��                          A                       5�_�                           ����                                                                                                                                                                                                                                                                                                                            %          +          V   #    f     �                         STOP_BITS : natural := 15��                          A       !               5�_�                            ����                                                                                                                                                                                                                                                                                                                            $          *          V   #    f     �                 5��                          A                      5�_�                           ����                                                                                                                                                                                                                                                                                                                            #          )          V   #    f     �         �              WIDTH: natural := 7 ;5��                        =                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            #          )          V   #    f     �         �              WIDTH: natural := 75��                         =                      �                        <                     �                         >                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f4     �         �      (        init: in bit_vector(7 downto 0);�         �    5��                        �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       f8     �      	   �      %        d: in bit_vector(7 downto 0);�      	   �    5��                        �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        fV     �                )    signal value: bit_vector(7 downto 0);�      
          %        q: out bit_vector(7 downto 0)�      	   �      %        d: in bit_vector(7 downto 0);5��                        �                     �                        �                     �                        _                    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        fe     �                .        init: in bit_vector(WIDTH-1 downto 0);5��                          s       /               5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        fq     �         �                  value <= init;5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        fu     �         �                  value <= ;5��                         �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        fu    �         �                  value <= ();5��                         �                     �                        �                    �                        �                    �                        �                    �                        �                    5�_�                       	    ����                                                                                                                                                                                                                                                                                                                                                  V        f�     �          �      use IEEE.STD_LOGIC_1164.ALL;5��       	                 x                    �       	                 x                    �       	                 x                    �       	                 x                    �       	                 x                    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        f�     �         �    5��                          M                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        f�     �      <   �    �         �    5��                          N              �      5�_�                             ����                                                                                                                                                                                                                                                                                                                                       )          V       f�     �   '   )          #architecture rtl of counter_6bit is�   %   '          end counter_6bit;�      !   �      entity counter_6bit is5��                        �                    �    %                    Y                    �    '                                        5�_�                     2       ����                                                                                                                                                                                                                                                                                                                            2          2   %       v   %    f=     �   1   3   �      +        elsif to_integer(counter) = 63 then�   2   3   �    5��    1                    T                    5�_�      !              3       ����                                                                                                                                                                                                                                                                                                                            2          2          v   %    fF     �   3   5   �    5��    3                      �                     �    3                      �                     5�_�       "           !   4        ����                                                                                                                                                                                                                                                                                                                            2          2          v   %    fF     �   3   5   �       �   4   5   �    5��    3                      �                     5�_�   !   #           "   5   
    ����                                                                                                                                                                                                                                                                                                                            2          2          v   %    fL     �   4   6   �      #        elsif rising_edge(clk) then5��    4                     �                     5�_�   "   $           #   5   	    ����                                                                                                                                                                                                                                                                                                                            2          2          v   %    fM     �   4   6   �      !        sif rising_edge(clk) then5��    4                    �                    5�_�   #   %           $   4        ����                                                                                                                                                                                                                                                                                                                            4           4          v       fV     �   3   5   �      to_integer(counter) = 635��    3                      �                     5�_�   $   &           %   5       ����                                                                                                                                                                                                                                                                                                                            5          5          v       fZ     �   4   6   �      $            if rising_edge(clk) then�   5   6   �    5��    4                    �                    5�_�   %   '           &   4        ����                                                                                                                                                                                                                                                                                                                            5          5   &       v       f[     �   3   4           5��    3                      �                     5�_�   &   (           '   5       ����                                                                                                                                                                                                                                                                                                                            4          4   &       v       f^     �   4   6   �      #            counter <= counter + 1;5��    4                     �                     5�_�   '   )           (   5       ����                                                                                                                                                                                                                                                                                                                            4          4   &       v       f_     �   5   8   �                      �   5   7   �    5��    5                      �                     �    5                     �                     �    5                     �                    �    5                    �                     �    6                     �                    5�_�   (   *           )   7       ����                                                                                                                                                                                                                                                                                                                            4          4   &       v       fm     �   6   7                          done5��    6                      �                     5�_�   )   +           *   5       ����                                                                                                                                                                                                                                                                                                                            4          4   &       v       fn     �   4   5          '                counter <= counter + 1;5��    4                      �      (               5�_�   *   -           +   5       ����                                                                                                                                                                                                                                                                                                                            4          4   &       v       fn     �   5   7   �    �   5   6   �    5��    5                      �              (       5�_�   +   .   ,       -   3       ����                                                                                                                                                                                                                                                                                                                            4          4   &       v       fs     �   2   3                      done <= '1';5��    2                      j                     5�_�   -   /           .   3       ����                                                                                                                                                                                                                                                                                                                            3          3   &       v       fs     �   3   5   �    �   3   4   �    5��    3                      �                     5�_�   .   0           /   4       ����                                                                                                                                                                                                                                                                                                                            3          3   &       v       ft     �   3   5   �                  done <= '1';5��    3                     �                     5�_�   /   2           0   6       ����                                                                                                                                                                                                                                                                                                                            3          3   &       v       fv     �   6   8   �                      �   6   8   �    5��    6                      �                     �    6                     �                     �    6                     �                    �    6                     �                     5�_�   0   3   1       2   3   '    ����                                                                                                                                                                                                                                                                                                                            3          3   &       v       f�     �   2   4   �      ,            if to_integer(counter) = 63 then5��    2   &                  �                     �    2   %                  �                     5�_�   2   4           3   3   %    ����                                                                                                                                                                                                                                                                                                                            3          3   &       v       f�     �   2   4   �      *            if to_integer(counter) =  then5��    2   %                  �                     5�_�   3   5           4   3   &    ����                                                                                                                                                                                                                                                                                                                            3          3   &       v       f�     �   2   4   �      ,            if to_integer(counter) = () then5��    2   &                  �                     �    2   &                 �                    �    2   &                 �                    �    2   &                 �                    �    2   &                 �                    5�_�   4   6           5   3   2    ����                                                                                                                                                                                                                                                                                                                            3          3   &       v       f�     �   2   4   �      9            if to_integer(counter) = (others => '0') then5��    2   1                 �                    5�_�   5   7           6   3       ����                                                                                                                                                                                                                                                                                                                            3          3   &       v       f�     �   2   4   �      9            if to_integer(counter) = (others => '1') then5��    2          
           y      
               5�_�   6   8           7   3       ����                                                                                                                                                                                                                                                                                                                            3          3   &       v       f�     �   2   4   �      /            if (counter) = (others => '1') then5��    2                     y                     5�_�   7   9           8   3       ����                                                                                                                                                                                                                                                                                                                            3          3   &       v       f�     �   2   4   �      .            if counter) = (others => '1') then5��    2                     �                     5�_�   8   :           9            ����                                                                                                                                                                                                                                                                                                                                                V       f�     �       $   �    �       !   �    5��                           �              0       5�_�   9   ;           :   '       ����                                                                                                                                                                                                                                                                                                                                                V       f     �   &   (   �      O        count : out unsigned(5 downto 0)       -- 6-bit count output (64 steps)5��    &                    ;                    5�_�   :   <           ;   ,       ����                                                                                                                                                                                                                                                                                                                                                V       f     �   +   -   �      )    signal counter: unsigned(5 downto 0);5��    +                     �                     5�_�   ;   =           <   ,       ����                                                                                                                                                                                                                                                                                                                                                V       f     �   +   -   �          signal counter: );5��    +                    �                    �    +                    �                    �    +                    �                    �    +                    �                    5�_�   <   >           =   6       ����                                                                                                                                                                                                                                                                                                                            6          6   '       v   '    f+     �   5   7   �      -            if counter = (others => '1') then5��    5                    �                    �    5                    �                    �    5                     �                     �    5                    �                    �    5                     �                     �    5                    �                    �    5                    �                    �    5                    �                    5�_�   =   ?           >   3       ����                                                                                                                                                                                                                                                                                                                            6          6   '       v   '    f5     �   2   4   �      '            counter <= (others => '0');5��    2                    2                    5�_�   >   @           ?   �        ����                                                                                                                                                                                                                                                                                                                            C          �           V       fO     �   B           l   library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity serial_out is       generic(   #        POLARITY : boolean := TRUE;           WIDTH: natural := 7 ;           PARITY : natural := 1 ;            STOP_BITS : natural := 1           );   	    port(   #        clk, reset, tx_go : in bit;           tx_done : out bit;   /        data : in bit_vector(WIDTH-1 downto 0);           serial_o : out bit       );   end serial_out;       (architecture Behavioral of serial_out is       type state_t is (           INICIO, START_BIT,   i        TRANSMISSAO0, TRANSMISSAO1, TRANSMISSAO2, TRANSMISSAO3, TRANSMISSAO4, TRANSMISSAO5, TRANSMISSAO6,           STOP_BIT   
        );   +    signal estado_atual: state_t := INICIO;   ,    signal prox_estado: state_t:= START_BIT;   "    signal enviados: integer := 0;           p1: process(clk) begin   "        if (rising_edge(clk)) then   (            estado_atual <= prox_estado;           end if;               if (reset = '1') then   #            estado_atual <= INICIO;   "            prox_estado <= INICIO;               enviados <= 0;           end if;               case estado_atual is                when INICIO =>                   tx_done <= '0';                    serial_o <= '1';                   enviados <= 0;   #                if tx_go = '1' then   -                    prox_estado <= START_BIT;                   else       *                    prox_estado <= INICIO;                   end if;                   when START_BIT =>                   tx_done <= '0';                    serial_o <= '0';   ,                prox_estado <= TRANSMISSAO0;                               when TRANSMISSAO0 =>                   tx_done <= '0';   $                serial_o <= data(0);   ,                prox_estado <= TRANSMISSAO1;                               when TRANSMISSAO1 =>                   tx_done <= '0';   $                serial_o <= data(1);   ,                prox_estado <= TRANSMISSAO2;                               when TRANSMISSAO2 =>                   tx_done <= '0';   $                serial_o <= data(2);   ,                prox_estado <= TRANSMISSAO3;                               when TRANSMISSAO3 =>                   tx_done <= '0';   $                serial_o <= data(3);   ,                prox_estado <= TRANSMISSAO4;                    when TRANSMISSAO4 =>                   tx_done <= '0';   $                serial_o <= data(4);   ,                prox_estado <= TRANSMISSAO5;                    when TRANSMISSAO5 =>                   tx_done <= '0';   $                serial_o <= data(5);   ,                prox_estado <= TRANSMISSAO6;                    when TRANSMISSAO6 =>                   tx_done <= '0';   $                serial_o <= data(6);   (                prox_estado <= STOP_BIT;                              when STOP_BIT =>                   tx_done <= '1';                    serial_o <= '1';   &                prox_estado <= INICIO;                   when others =>   &                prox_estado <= INICIO;               end case;       end process p1;   end architecture;                            5��    B       l       l       r            >      5�_�   ?   A           @   �        ����                                                                                                                                                                                                                                                                                                                            C          �           V       fR    �   �   �          --   --   --   --   --   --5��    �                      �                     5�_�   @   B           A           ����                                                                                                                                                                                                                                                                                                                            C          �           V       f�    �          �    �         �    5��                                           )       5�_�   A   C           B   �       ����                                                                                                                                                                                                                                                                                                                            F          �          V       f     �   E           f   -- library IEEE;   -- use IEEE.NUMERIC_BIT.ALL;   --   -- entity serial_out is   --     generic(   &--         POLARITY : boolean := TRUE;    --         WIDTH: natural := 7 ;   "--         PARITY : natural := 1 ;   #--         STOP_BITS : natural := 1   --   	--     );   --     port(   &--         clk, reset, tx_go : in bit;   --         tx_done : out bit;   2--         data : in bit_vector(WIDTH-1 downto 0);   --         serial_o : out bit   	--     );   -- end serial_out;   --   +-- architecture Behavioral of serial_out is   --     type state_t is (   --         INICIO, START_BIT,   l--         TRANSMISSAO0, TRANSMISSAO1, TRANSMISSAO2, TRANSMISSAO3, TRANSMISSAO4, TRANSMISSAO5, TRANSMISSAO6,   --         STOP_BIT   --         );   .--     signal estado_atual: state_t := INICIO;   /--     signal prox_estado: state_t:= START_BIT;   %--     signal enviados: integer := 0;   --   --     p1: process(clk) begin   %--         if (rising_edge(clk)) then   +--             estado_atual <= prox_estado;   --         end if;   --    --         if (reset = '1') then   &--             estado_atual <= INICIO;   %--             prox_estado <= INICIO;   --             enviados <= 0;   --         end if;   --    --         case estado_atual is    --             when INICIO =>   "--                 tx_done <= '0';   #--                 serial_o <= '1';   !--                 enviados <= 0;   &--                 if tx_go = '1' then   0--                     prox_estado <= START_BIT;   --                 else       ---                     prox_estado <= INICIO;   --                 end if;   --    --             when START_BIT =>   "--                 tx_done <= '0';   #--                 serial_o <= '0';   /--                 prox_estado <= TRANSMISSAO0;   --                #--             when TRANSMISSAO0 =>   "--                 tx_done <= '0';   '--                 serial_o <= data(0);   /--                 prox_estado <= TRANSMISSAO1;   --                #--             when TRANSMISSAO1 =>   "--                 tx_done <= '0';   '--                 serial_o <= data(1);   /--                 prox_estado <= TRANSMISSAO2;   --                #--             when TRANSMISSAO2 =>   "--                 tx_done <= '0';   '--                 serial_o <= data(2);   /--                 prox_estado <= TRANSMISSAO3;   --                #--             when TRANSMISSAO3 =>   "--                 tx_done <= '0';   '--                 serial_o <= data(3);   /--                 prox_estado <= TRANSMISSAO4;   --   #--             when TRANSMISSAO4 =>   "--                 tx_done <= '0';   '--                 serial_o <= data(4);   /--                 prox_estado <= TRANSMISSAO5;   --   #--             when TRANSMISSAO5 =>   "--                 tx_done <= '0';   '--                 serial_o <= data(5);   /--                 prox_estado <= TRANSMISSAO6;   --   #--             when TRANSMISSAO6 =>   "--                 tx_done <= '0';   '--                 serial_o <= data(6);   +--                 prox_estado <= STOP_BIT;   --                --             when STOP_BIT =>   "--                 tx_done <= '1';   #--                 serial_o <= '1';   )--                 prox_estado <= INICIO;   --   --             when others =>   )--                 prox_estado <= INICIO;   --             end case;   --     end process p1;   -- end architecture;   --5��    E       f       f       �      ,            5�_�   B   D           C   X        ����                                                                                                                                                                                                                                                                                                                            F          �          V       f*�     �   ^   `   �      end architecture �   X   Z   �      architecture rtl of  is�   \   `   �          �   X   ^   �      arch�   W   Z   �       �   W   Y   �    5��    W                                           �    W                                           �    X                                           �    X                                          �    X                                          �    X                                         �    X                                         �    X                                         �    X                                         �    X                    1                     �    \                      I                      �    \                    I                     �    ^                     `                     �    X                     1                     �    ^                     k                     5�_�   C   E           D   Y       ����                                                                                                                                                                                                                                                                                                                            Y          Y          v       f*�     �   Y   Z   �    �   ^   `   �      end architecture rtl;�   X   Z   �      "architecture rtl of transmissao is�   Y   Z   �    �   Y   Z   �    �   Y   Z   �    �   Y   Z   �    �   Y   Z   �    �   Y   Z   �    �   Y   Z   �    5��    X                    *                    �    ^                    i                    �    X                     +                     �    ^                    j                    �    X                     ,                     �    ^                    k                    �    X                     -                     �    ^                    l                    �    X                     -                     �    ^                    k                    �    X                     ,                     �    ^                    j                    �    X                     +                     �    ^                    i                    �    X                 
   *             
       �    X          
          *      
              �    X                 
   *             
       �    ^                 
   r             
       5�_�   D   F           E   Y       ����                                                                                                                                                                                                                                                                                                                            Y   %       Y          v       f+     �   \   ^   �          �   X   Z   �      )architecture Behavioral of transmissao is5��    X                    8                    �    X                     :                     �    X                     9                     �    X                 
   8             
       �    X          
          8      
              �    X                 
   8             
       �    \                     Z                     5�_�   E   G           F   Z       ����                                                                                                                                                                                                                                                                                                                            Y   %       Y          v       f+     �   Y   \   �          �   Y   [   �    5��    Y                      F                     �    Y                      F                     �    Y                     F                     �    Z                  	   K              	       �    Z                    S                    5�_�   F   H           G   [       ����                                                                                                                                                                                                                                                                                                                            Y   %       Y          v       f+-     �   Z   \   �          component �   [   \   �    5��    Z                     U                     5�_�   G   I           H   [       ����                                                                                                                                                                                                                                                                                                                            Y   %       Y          v       f+.     �   Z   ]   �          component generic_reg5��    Z                     `                     �    Z                    c                     �    [                     d                    �    [                      d                     5�_�   H   J           I   [        ����                                                                                                                                                                                                                                                                                                                                                  V        f+�     �   [   d   �    �   [   \   �    5��    [                      d              �       5�_�   I   K           J   \       ����                                                                                                                                                                                                                                                                                                                            \          c                 f+�     �   \   d   �              WIDTH: natural := 8       );   
    port (   !        rst, clk, enable: in bit;   +        d: in bit_vector(WIDTH-1 downto 0);   +        q: out bit_vector(WIDTH-1 downto 0)       );�   [   ]   �          generic(5��    [                     h                     �    \                     y                     �    ]                     �                     �    ^                     �                     �    _                     �                     �    `                     �                     �    a                     	                     �    b                     9                     5�_�   J   M           K   d        ����                                                                                                                                                                                                                                                                                                                            \          c                 f+�     �   c   e   �       5��    c                      @                     �    c                     @                    �    c                     H                     �    c   
                  J                     �    c   	                  I                     �    c                 	   H             	       �    c          	          H      	              �    c                 
   H             
       5�_�   K   N   L       M   [       ����                                                                                                                                                                                                                                                                                                                            \          c                 f+�     �   Z   \   �          component generic_reg is5��    Z                     `                     5�_�   M   O           N   d       ����                                                                                                                                                                                                                                                                                                                            d          [          V       f+�     �   d   f   �    5��    d                      P                     �    d                      P                     5�_�   N   P           O   e        ����                                                                                                                                                                                                                                                                                                                            d          [          V       f+�     �   e   p   �    �   e   f   �    5��    e               
       Q              	      5�_�   O   Q           P   f       ����                                                                                                                                                                                                                                                                                                                            d          [          V       f+�     �   e   g   �          component generic_reg5��    e                    _                    �    e                    _                    �    e                    _                    �    e                    _                    �    e                    _                    5�_�   P   R           Q   g        ����                                                                                                                                                                                                                                                                                                                            g          n   
       V       f+�     �   f   o   �    �   g   h   �    �   f   g                  generic(               WIDTH: natural := 8   
        );           port (   %            rst, clk, enable: in bit;   /            d: in bit_vector(WIDTH-1 downto 0);   /            q: out bit_vector(WIDTH-1 downto 0)   
        );5��    f                      o      �               �    f                      o              �       5�_�   Q   S           R   g       ����                                                                                                                                                                                                                                                                                                                            g          n                 f+�     �   g   o   �              WIDTH: natural := 8       );   
    port (   C        clk, rst: in bit;                            -- Clock input           done: out bit;   B        count : out natural       -- 6-bit count output (64 steps)       );�   f   h   �          generic(5��    f                     s                     �    g                     �                     �    h                     �                     �    i                     �                     �    j                     �                     �    k                     	                     �    l                     !	                     �    m                     h	                     5�_�   R   T           S   ]       ����                                                                                                                                                                                                                                                                                                                            g          n                 f,<     �   \   ^   �                  WIDTH: natural := 85��    \                     �                     �    \                     �                     �    \                     �                     �    \                     �                     5�_�   S   U           T   h       ����                                                                                                                                                                                                                                                                                                                            g          n                 f,J     �   g   i   �                  WIDTH: natural := 85��    g                     �                     �    g                     �                     �    g                     �                     �    g                     �                     5�_�   T   V           U   %       ����                                                                                                                                                                                                                                                                                                                            g          n                 f,R     �   $   &   �              WIDTH: natural := 85��    $                     �                     �    $                     �                     �    $                     �                     �    $                     �                     �    $                     �                     5�_�   U   W           V   %       ����                                                                                                                                                                                                                                                                                                                            g          n                 f,W     �   $   &   �              WIDTH: natural5��    $                    �                    �    $                     �                     5�_�   V   X           W   9       ����                                                                                                                                                                                                                                                                                                                            9          9          v       f,e    �   8   :   �      %            if counter = WIDTH-1 then�   9   :   �    5��    8                 	   �             	       5�_�   W   Y           X   L       ����                                                                                                                                                                                                                                                                                                                            9          9   !       v       f,�     �   K   M   �              WIDTH: natural := 7 ;5��    K                     (                     5�_�   X   Z           Y   M       ����                                                                                                                                                                                                                                                                                                                            9          9   !       v       f,�     �   L   N   �              PARITY : natural := 1 ;5��    L                     G                     5�_�   Y   \           Z   O        ����                                                                                                                                                                                                                                                                                                                            9          9   !       v       f,�     �   N   O           5��    N                      j                     5�_�   Z   ]   [       \   n       ����                                                                                                                                                                                                                                                                                                                            9          9   !       v       f-     �   o   q   �      
    signal�   n   q   �          �   n   p   �    5��    n                      x	                     �    n                      x	                     �    n                     x	                     �    o                     }	                     �    o                     �	                     �    o                     	                     �    o                     ~	                     �    o                    }	                    �    o                    }	                    �    o                    }	                    5�_�   \   ^           ]   p       ����                                                                                                                                                                                                                                                                                                                            9          9   !       v       f-     �   o   q   �          signal i: natural;5��    o                    �	                    �    o                     �	                     5�_�   ]   _           ^   t       ����                                                                                                                                                                                                                                                                                                                            9          9   !       v       f-     �   s   u   �          kj5��    s                     �	                     �    s                     �	                     �    s                     �	                     �    s                     �	                     �    s                      �	                     5�_�   ^   `           _   p       ����                                                                                                                                                                                                                                                                                                                            9          9   !       v       f->     �   p   r   �          �   p   r   �    5��    p                      �	                     �    p                     �	                     �    p                    �	                    5�_�   _   a           `   u        ����                                                                                                                                                                                                                                                                                                                            9          9   !       v       f-N     �   u   x   �              �   t   w   �       5��    t                      �	                     �    t                     �	                     �    t                    �	                    �    t                     �	                     �    t                    �	                    �    t                    �	                    �    t                    �	                    �    t                    �	                    �    t                    �	                     �    u                      �	                      �    u                    �	                     5�_�   `   b           a   u       ����                                                                                                                                                                                                                                                                                                                            u          u          v       f-h     �   t   v   �          if condition then5��    t          	          �	      	              5�_�   a   c           b   v        ����                                                                                                                                                                                                                                                                                                                            u   	       w   	       V   	    f-�     �   w   y   �          end process �   v   y   �              �   t   x   �          if rst then�   u   v                         end if;5��    u                      �	                     �    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t   
                  �	                     �    t   	                  �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t   
                  �	                     �    t   	                  �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t   
                  �	                     �    t   	                  �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t   
                  �	                     �    t   	                  �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t   
                  �	                     �    t   	                  �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t   
                  �	                     �    t   	                  �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t   
                  �	                     �    t   	                  �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t   
                  �	                     �    t   	                  �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t   
                  �	                     �    t   	                  �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t   
                  �	                     �    t   	                  �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t   
                  �	                     �    t   	                  �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t   
                  �	                     �    t   	                  �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                    �	                    �    t                    �	                    �    t                 #   �	             #       �    t   '                 �	                     �    v                      �	                      �    v                    �	                     �    w                  
   
              
       5�_�   b   d           c   u       ����                                                                                                                                                                                                                                                                                                                            u          u          v       f-�     �   w   y   �          end process proc_name;�   t   v   �      (    proc_name: process(sensitivity_list)5��    t          	           �	      	               �    w          	           �	      	               5�_�   c   e           d   u       ����                                                                                                                                                                                                                                                                                                                            u          u          v       f-�     �   t   v   �          : process(sensitivity_list)5��    t                     �	                     5�_�   d   f           e   u       ����                                                                                                                                                                                                                                                                                                                            u          u          v       f-�     �   t   v   �          process(sensitivity_list)5��    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                    �	                    �    t                    �	                    �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                     �	                     �    t                    �	                    �    t                    �	                    �    t                    �	                    5�_�   e   g           f   u        ����                                                                                                                                                                                                                                                                                                                            u          u          v       f-�     �   t   u              process(reset)   	    begin           5��    t                      �	      &               5�_�   f   h           g   u        ����                                                                                                                                                                                                                                                                                                                            u          u          v       f-�    �   t   u              end process ;       5��    t                      �	                     5�_�   g   i           h   s        ����                                                                                                                                                                                                                                                                                                                                                             f/�     �   u   w   �              generic�   s   w   �          �   s   u   �    5��    s                      �	                     �    s                      �	                     �    s                      �	                     �    s                     �	                     �    t                  	   �	              	       �    t                     �	                     �    t                    �	                     �    u                     �	                     �    u   
                  �	                     �    u   	                  �	                     �    u                    �	                    �    u   
                  �	                     �    u   	                  �	                     �    u                    �	                    �    u                    �	                    �    u                    �	                    5�_�   h   j           i   v       ����                                                                                                                                                                                                                                                                                                                                                             f/�     �   u   w   �              generic map5��    u                     �	                     5�_�   i   k           j   u       ����                                                                                                                                                                                                                                                                                                                                                             f/�     �   t   v   �          counter:5��    t                     �	                     �    t                    �	                    �    t                    �	                    �    t                    �	                    �    t                    �	                    �    t                    �	                    �    t                    �	                    �    t                    �	                    5�_�   j   l           k   v       ����                                                                                                                                                                                                                                                                                                                                                             f/�     �   u   w   �              generic map()5��    u                     �	                     �    u                    �	                    �    u                    �	                    �    u                    �	                    5�_�   k   m           l   v       ����                                                                                                                                                                                                                                                                                                                                                             f/�     �   v   x   �              port�   u   x   �              generic map(WIDTH)5��    u                     �	                     �    u                    �	              	       �    v                     �	                     �    v   
                  �	                     �    v   	                  �	                     �    v                    �	                    �    v                    �	                    �    v                    �	                    5�_�   l   n           m   g       ����                                                                                                                                                                                                                                                                                                                                                             f/�     �   f   h   �                  WIDTH: natural5��    f                    �                    �    f                 	   �             	       �    f          	       	   �      	       	       �    f          	          �      	              �    f                 	   �             	       5�_�   m   o           n   w       ����                                                                                                                                                                                                                                                                                                                                                             f/�     �   v   x   �              port map5��    v                     �	                     5�_�   n   p           o   v       ����                                                                                                                                                                                                                                                                                                                                                             f/�     �   u   w   �              generic map(WIDTH);5��    u                     �	                     5�_�   o   q           p   w       ����                                                                                                                                                                                                                                                                                                                                                             f/�     �   v   x   �              port map()5��    v                     �	                     �    v                     
                     �    v                     
                     �    v                    
                    �    v                    �	                    �    v                    �	                    �    v                    �	                    �    v                     �	                     5�_�   p   r           q   Q       ����                                                                                                                                                                                                                                                                                                                                                             f0     �   P   R   �      #        clk, reset, tx_go : in bit;5��    P                    �                    5�_�   q   s           r   j   <    ����                                                                                                                                                                                                                                                                                                                                                             f0     �   i   k   �      G            clk, rst: in bit;                            -- Clock input5��    i   <                 �                    5�_�   r   t           s   w       ����                                                                                                                                                                                                                                                                                                                                                             f00     �   v   x   �              port map()5��    v                     
                     5�_�   s   u           t   w   '    ����                                                                                                                                                                                                                                                                                                                                                             f0=     �   v   x   �      '        port map(clock, reset, done, i)5��    v   '                  
                     5�_�   t   v           u   u       ����                                                                                                                                                                                                                                                                                                                                                             f0G     �   t   v   �          counter: counter_generic5��    t                    �	                    �    t                    �	                    5�_�   u   w           v   v       ����                                                                                                                                                                                                                                                                                                                                                             f0�     �   u   w   �              generic map(WIDTH)5��    u                     �	                     5�_�   v   x           w   w       ����                                                                                                                                                                                                                                                                                                                                                             f2S     �   {   }   �          end process �   z   }   �              �   x   |   �          cproc, processc�   w   z   �              �   w   y   �    5��    w                       
              	       �    w                       
                     �    w                      
              	       �    x                    %
                    �    x                    &
                    �    x                    &
                    �    x                     &
                     �    x                    %
                    �    x                     &
                     �    x                    %
                    �    x                     ,
                     �    x   
                  +
                     �    x   	                  *
                     �    x                     )
                     �    x                     (
                     �    x                     '
                     �    x                     &
                     �    x                    %
                    �    x                    %
                    �    x                    %
                    �    x                 #   %
             #       �    x   '                 H
                     �    z                      \
                      �    z                    \
                     �    {                  
   m
              
       5�_�   w   y           x   y       ����                                                                                                                                                                                                                                                                                                                            y          y          v       f2o     �   y   z   �    �   {   }   �          end process proc_name;�   y   z   �    �   y   z   �    �   y   z   �    �   y   z   �    �   y   z   �    �   y   z   �    �   y   z   �    �   y   z   �    �   y   z   �    �   y   z   �    �   y   z   �    �   y   z   �    �   y   z   �    �   y   z   �    �   y   z   �    �   y   z   �    �   x   z   �      (    proc_name: process(sensitivity_list)5��    x          	          %
      	              �    {          	          e
      	              �    x                     &
                     �    {                    f
                    �    x                     &
                     �    x                    %
                    �    {                    g
                    �    x                     '
                     �    x                     &
                     �    x                    %
                    �    {                    h
                    �    x                     (
                     �    x                     '
                     �    x                     &
                     �    x                    %
                    �    {                    k
                    �    x   
                  +
                     �    x   	                  *
                     �    x                     )
                     �    x                     (
                     �    x                     '
                     �    x                     &
                     �    x                 	   %
             	       �    {                 	   m
             	       �    x                     -
                     �    {          	          l
      	              �    x                     ,
                     �    {                    k
                    �    x   
                  +
                     �    {                    j
                    �    x   	                  *
                     �    {                    i
                    �    x                     )
                     �    {                    h
                    �    x                     (
                     �    {                    g
                    �    x                     '
                     �    {                    f
                    �    x                     &
                     �    {                    e
                    �    x                     %
                     �    {                     d
                     �    x                     %
                     �    {                     e
                     �    x                     &
                     �    {                    f
                    5�_�   x   z           y   y       ����                                                                                                                                                                                                                                                                                                                            y          y          v       f2z     �   {   ~   �                  �   z   }   �              �   x   z   �      !    lg: process(sensitivity_list)5��    x                    1
                    �    x                     3
                     �    x                    2
                    �    x                     <
                     �    x                     ;
                     �    x                     :
                     �    x                     9
                     �    x                    8
                    �    x                    8
                    �    x                    8
                    �    z                     Q
                     �    z   	                  R
                     �    z                    Q
                    �    z   	                  R
                     �    z                    Q
                    �    z                    Q
                    �    z                    Q
                    �    z                    Q
                    �    z                    ]
                     �    {                      o
                      �    {                    o
                     5�_�   y   {           z   {       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f2�     �   z   |   �              if condition then5��    z          	          T
      	              �    z                     V
                     �    z                     U
                     �    z                    T
                    �    z                    T
                    �    z                 	   T
             	       �    z                     \
                     5�_�   z   |           {   {       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f2�     �   z   |   �              if reset =  then5��    z                     \
                     5�_�   {   }           |   {       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f2�     �   {   }   �                  done�   z   |   �              if reset = '' then5��    z                     ]
                     �    {                     q
                     �    {                    r
                    �    {                     s
                     �    {                     r
                     �    {                    q
                    �    {                    q
                    �    {                    q
                    5�_�   |   ~           }   |       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f2�     �   {   }   �                  done <= 5��    {                     y
                     5�_�   }              ~   |       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f2�     �   {   }   �                  done <= ''5��    {                     z
                     5�_�   ~   �              |       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f2�     �   |   ~   �                  tx_done�   {   ~   �                  done <= '1'5��    {                     |
                     �    {                    }
                     �    |                     �
                     �    |                     �
                     �    |                    �
                    �    |                     �
                     �    |                     �
                     �    |                     �
                     �    |                     �
                     �    |                     �
                     �    |                     �
                     �    |                    �
                    �    |                    �
                    �    |                    �
                    5�_�      �           �   }       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f2�     �   |   ~   �                  tx_done <= 5��    |                     �
                     5�_�   �   �           �   }       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f2�     �   |   ~   �                  tx_done <= ''5��    |                     �
                     5�_�   �   �           �   }       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f2�     �   |   ~   �                  tx_done <= '1'5��    |                     �
                     5�_�   �   �   �       �   v       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f2�     �   u   w   �              generic map(WIDTH+1)5��    u                     �	                     �    u                     �	                    �    u   ,                  
                     5�_�   �   �           �   v       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f2�     �   u   w   �      B    generic map(WIDTH+1)    -- The plus 1 is to send the start bit5��    u                     �	                     5�_�   �   �           �   v       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3P     �   u   w   �      F        generic map(WIDTH+1)    -- The plus 1 is to send the start bit5��    u                     �	                     5�_�   �   �           �   v       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3a     �   u   w   �      G        generic map(WIDTH+1+)    -- The plus 1 is to send the start bit�   v   w   �    5��    u                  	   �	              	       5�_�   �   �           �   v   P    ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3d     �   u   w   �      P        generic map(WIDTH+1+STOP_BITS)    -- The plus 1 is to send the start bit5��    u   M                 '
                    5�_�   �   �           �   v   7    ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3j     �   u   w   �      Z        generic map(WIDTH+1+STOP_BITS)    -- The plus 1 is to send the start and stop bits5��    u   5                 
                    �    u   5                  
                     5�_�   �   �           �   v   5    ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3o     �   u   w   �      X        generic map(WIDTH+1+STOP_BITS)    -- The plus is to send the start and stop bits5��    u   1                 
                    5�_�   �   �           �   v   6    ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3u     �   u   w   �      X        generic map(WIDTH+1+STOP_BITS)    -- The sums is to send the start and stop bits5��    u   6                 
                    5�_�   �   �           �   v   L    ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3�     �   u   w   �      Y        generic map(WIDTH+1+STOP_BITS)    -- The sums are to send the start and stop bits5��    u   K                 %
                    5�_�   �   �           �   v   M    ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3�     �   u   w   �      V        generic map(WIDTH+1+STOP_BITS)    -- The sums are to send the start, stop bits5��    u   M                  '
                     5�_�   �   �           �   v       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3�     �   u   w   �      a        generic map(WIDTH+1+STOP_BITS)    -- The sums are to send the start, parity and stop bits5��    u                    �	                    5�_�   �   �           �   }       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3�     �   }      �                  �   }      �    5��    }                      �
                     �    }                     �
                     �    }                     �
                     �    }                     �
                     �    }                    �
                    �    }                    �
                    �    }                     �
                     �    }                     �
                     �    }                     �
                     �    }                     �
                     �    }                    �
                    �    }                    �
                    �    }                    �
                    5�_�   �   �           �   ~       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3�     �   }      �                  elsif5��    }                     �
                     5�_�   �   �           �   ~       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3�     �   }      �              elsif5��    }                     �
                     �    }                     �
                     �    }                     �
                     �    }                    �
                    �    }                    �
                    �    }                    �
                    5�_�   �   �           �   ~       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3�     �   }      �              elsif rising_edge5��    }                     �
                     5�_�   �   �           �   ~       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3�     �   }      �              elsif rising_edge()5��    }                     �
                     �    }                    �
                    �    }                    �
                    �    }                    �
                    5�_�   �   �           �   ~        ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3�     �   }      �               elsif rising_edge(clock)5��    }                      �
                     5�_�   �   �           �   ~   %    ����                                                                                                                                                                                                                                                                                                                            {          {          v       f3�     �   ~   �   �                  if tx_done�   }   �   �      %        elsif rising_edge(clock) then5��    }   %                               	       �    ~                                         �    ~                                          �    ~                                          �    ~                                          �    ~                                          �    ~                                        �    ~                                          �    ~                                        �    ~                                        �    ~                                        �    ~                                          �    ~                                          �    ~                                          �    ~                                        �    ~                                          �    ~                                          �    ~                                          �    ~                                          �    ~                                        �    ~                                        �    ~                                        �    ~                                          �    ~                                          5�_�   �   �           �   q       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f4�     �   p   r   �          signal done: bit;5��    p                    �	                    5�_�   �   �           �   w       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f4�     �   v   x   �      (        port map(clock, reset, done, i);5��    v                    ]
                    5�_�   �   �           �   w   %    ����                                                                                                                                                                                                                                                                                                                            {          {          v       f4�     �   v   x   �      *        port map(clock, reset, finish, i);5��    v   %                  c
                     5�_�   �   �           �   q       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f4�     �   p   r   �          signal finish: bit;5��    p                     �	                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            {          {          v       f4�     �   ~   �   �                  if tx_go and 5��    ~                     &                     �    ~                     )                     �    ~                     (                     �    ~                     '                     �    ~                    &                    �    ~                    &                    �    ~                    &                    �    ~   "                 /                    �    ~   "                 /                    �    ~   "                 /                    �    ~   &                 3                     �                         4                    �                          4                     �    ~   &                  3                     �    ~   %                  2                     �    ~   $                  1                     �    ~   #                  0                     �    ~   "                  /                     �    ~   !                  .                     �    ~                      -                     �    ~                     ,                     �    ~                     +                     �    ~                     *                     �    ~                     )                     �    ~                     (                     �    ~                     '                     �    ~                     &                     5�_�   �   �           �   q       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f5     �   p   q              signal finished: bit;5��    p                      �	                     5�_�   �   �           �   v       ����                                                                                                                                                                                                                                                                                                                            z          z          v       f5     �   u   w   �      ,        port map(clock, reset, finished, i);5��    u                    E
                    �    u                    E
                    �    u                    E
                    �    u                    E
                    �    u                    E
                    �    u                    E
                    5�_�   �   �           �   p       ����                                                                                                                                                                                                                                                                                                                            z          z          v       f8Q     �   p   r   �          �   p   r   �    5��    p                      �	                     �    p                     �	                     �    p                     �	                     �    p                    �	                    5�_�   �   �           �   w       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f8z     �   v   x   �      +        port map(clock, reset, tx_done, i);5��    v                    b
                    �    v   $                  g
                     �    v   #                 f
                    �    v   #                 f
                    �    v   #                 f
                    5�_�   �   �           �   j       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f95     �   i   k   �      G            clk, rst: in bit;                            -- clock input5��    i                     �                     5�_�   �   �           �   w       ����                                                                                                                                                                                                                                                                                                                            {          {          v       f9�     �   y   {   �              generic�   x   {   �          counting_state: generic_reg�   w   z   �              �   w   y   �    5��    w                      
              	       �    w                      
                     �    w                     
              	       �    x                    �
                    �    x                     �
                     �    x                     �
                     �    x                    �
                    �    x                     �
                     �    x                     �
                     �    x                     �
                     �    x                     �
                     �    x                     �
                     �    x                     �
                     �    x                    �
                    �    x                     �
                     �    x                     �
                     �    x                     �
                     �    x                     �
                     �    x                     �
                     �    x                     �
                     �    x                     �
                     �    x                     �
                     �    x                     �
                     �    x                     �
                     �    x                    �
                    �    x                    �
                    �    x                    �
                    �    x                    �
                     �    y                     �
                     �    y                    �
                    �    y                    �
                    �    y                     �
                     �    y                     �
                     �    y                     �
                     �    y                     �
                     �    y   
                  �
                     �    y   	                  �
                     �    y                    �
                    �    y                    �
                    �    y                 
   �
             
       �    y                    �
                    5�_�   �   �           �   z       ����                                                                                                                                                                                                                                                                                                                            ~          ~          v       f:-     �   y   {   �              generic map5��    y                     �
                     5�_�   �   �           �   z       ����                                                                                                                                                                                                                                                                                                                            ~          ~          v       f:1     �   y   {   �              generic map()5��    y                     �
                     5�_�   �   �           �   z       ����                                                                                                                                                                                                                                                                                                                            ~          ~          v       f:3     �   z   |   �              port�   y   |   �              generic map(1)5��    y                    �
              	       �    z                     �
                     �    z                    �
                    �    z                    �
                    �    z                    �
                    5�_�   �   �           �   {       ����                                                                                                                                                                                                                                                                                                                                                v       f:8     �   z   |   �              port map5��    z                     �
                     5�_�   �   �           �   {       ����                                                                                                                                                                                                                                                                                                                                                v       f:=     �   z   |   �              port map()5��    z                     �
                     �    z                    �
                    �    z                    �
                    �    z                    �
                    �    z                    �
                    �    z                    �
                    �    z                    �
                    �    z          	          �
      	              �    z                    �
                    �    z                    �
                    �    z                    �
                    �    z                 
   �
             
       �    z                    �
                    �    z                    �
                    �    z                 	   �
             	       �    z                      �
                     �    z                     �
                     5�_�   �   �           �   y       ����                                                                                                                                                                                                                                                                                                                            {          y          V       f˄     �   x   |   �          counting_state: generic_reg           generic map(1)            port map(reset, clock, )5��    x                     �
      X       a       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            {          y          V       fˉ     �   �   �   �                  if tx_go and 5��    �                    �                    �    �                     �                     �    �                    �                    �    �                     �                     �    �                 	   �             	       �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            {          y          V       f��     �   �   �   �                  �   �   �   �    5��    �                      [                     �    �                     g                     �    �                     h                     �    �                    g                    �    �                    g                    �    �                    g                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            {          y          V       f��     �   �   �   �                  is_counting <= 5��    �                     v                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            {          y          V       f��     �   �   �   �                  is_counting <= ''5��    �                     w                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            {          y          V       f��     �   �   �   �                  is_counting <= '0'5��    �                     y                     5�_�   �   �           �   �   $    ����                                                                                                                                                                                                                                                                                                                            {          y          V       f��     �   �   �   �      $            if i = 0 and is_counting5��    �   $                  �                     5�_�   �   �           �   �   '    ����                                                                                                                                                                                                                                                                                                                            {          y          V       f��     �   �   �   �      '            if i = 0 and is_counting = 5��    �   '                  �                     5�_�   �   �           �   �   (    ����                                                                                                                                                                                                                                                                                                                            {          y          V       f��     �   �   �   �      )            if i = 0 and is_counting = ''5��    �   (                  �                     5�_�   �   �           �   �   *    ����                                                                                                                                                                                                                                                                                                                            {          y          V       f��     �   �   �   �      *            if i = 0 and is_counting = '0'5��    �   *                  �                     �    �   +                 �                    �    �   +                 �                    �    �   +                 �                    �    �   /                 �                     �    �                     �                    �    �                      �                     5�_�   �   �           �   }       ����                                                                                                                                                                                                                                                                                                                            {          y          V       f�_     �   |   ~   �              �   |   ~   �    5��    |                      �
                     �    |                     �
                    �    |                    �
                    5�_�   �   �           �   }       ����                                                                                                                                                                                                                                                                                                                            {          y          V       f�f     �   |   ~   �          done <= 5��    |                     �
                     5�_�   �   �           �   }       ����                                                                                                                                                                                                                                                                                                                            {          y          V       f�f     �   |   ~   �          done <= ''5��    |                     �
                     5�_�   �   �           �   }       ����                                                                                                                                                                                                                                                                                                                            {          y          V       f�h     �   |   ~   �          done <= '1'5��    |                     �
                     �    |                     �
                    �    |                     �
                     �    |                     �
                     �    |                     �
                     �    |                     �
                     �    |                    �
                    �    |                    �
                    �    |                    �
                    5�_�   �   �           �   }   !    ����                                                                                                                                                                                                                                                                                                                            {          y          V       f�o     �   |   ~   �      !        done <= '1' when reset = 5��    |   !                                       5�_�   �   �           �   }   "    ����                                                                                                                                                                                                                                                                                                                            {          y          V       f�o     �   |   ~   �      #        done <= '1' when reset = ''5��    |   "                                       5�_�   �   �           �   }   $    ����                                                                                                                                                                                                                                                                                                                            {          y          V       f�p     �   |   ~   �      $        done <= '1' when reset = '1'5��    |   $                                       5�_�   �   �           �   }       ����                                                                                                                                                                                                                                                                                                                            {          y          V       f�r     �   |   ~   �      %        done <= '1' when reset = '1';5��    |                     �
                     �    |                     �
                     �    |                     �
                     �    |                     �
                     5�_�   �   �           �   q       ����                                                                                                                                                                                                                                                                                                                            {          y          V       fϙ     �   p   r   �          signal is_counting: bit;5��    p                    �	                    5�_�   �   �           �   j       ����                                                                                                                                                                                                                                                                                                                            {          y          V       f��     �   i   k   �      O            clk, rst, enable: in bit;                            -- clock input5��    i                    �                    5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                            {          y          V       f��     �   '   )   �      C        clk, rst: in bit;                            -- Clock input5��    '                                          5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            {          y          V       fЩ     �   /   1   �          �   /   1   �    5��    /                      �                     �    /                     �                     �    /                                          �    /                                          �    /                     
                     �    /                     	                     �    /                                          �    /                                          �    /                                          �    /                                        �    /                                          �    /                                        �    /                                        �    /                                        5�_�   �   �           �   8       ����                                                                                                                                                                                                                                                                                                                            |          z          V       fл     �   8   :   �                  �   8   :   �    5��    8                      �                     �    8                     �                     �    8                    �                    �    8                     �                     �    8                     �                     �    8                     �                     �    8                    �                    �    8                    �                    �    8                    �                    5�_�   �   �           �   9       ����                                                                                                                                                                                                                                                                                                                            }          {          V       f��     �   8   :   �                  is_counting <= 5��    8                     �                     5�_�   �   �           �   9       ����                                                                                                                                                                                                                                                                                                                            }          {          V       f��     �   8   :   �                  is_counting <= ''5��    8                     �                     5�_�   �   �           �   9       ����                                                                                                                                                                                                                                                                                                                            }          {          V       f��     �   8   :   �                  is_counting <= '0'5��    8                     �                     5�_�   �   �           �   =       ����                                                                                                                                                                                                                                                                                                                            }          {          V       f��     �   <   >   �                  else5��    <                    4                    �    <                    7                    �    <                     :                     �    <                     9                     �    <                     8                     �    <                    7                    �    <                    7                    �    <                    7                    5�_�   �   �           �   =        ����                                                                                                                                                                                                                                                                                                                            }          {          V       f��     �   <   >   �                   elsif is_counting = 5��    <                      E                     5�_�   �   �           �   =   !    ����                                                                                                                                                                                                                                                                                                                            }          {          V       f��     �   <   >   �      "            elsif is_counting = ''5��    <   !                  F                     5�_�   �   �           �   <       ����                                                                                                                                                                                                                                                                                                                            }          {          V       f��     �   <   >   �                      �   <   >   �    5��    <                      %                     �    <                     5                     �    <                     7                     �    <                     6                     �    <                    5                    �    <                    5                    �    <                    5                    �    <                     D                     5�_�   �   �           �   =       ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f��     �   <   >   �                      is_counting <= 5��    <                     D                     5�_�   �   �           �   =        ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f��     �   <   >   �      !                is_counting <= ''5��    <                      E                     5�_�   �   �           �   =   "    ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f��     �   <   >   �      "                is_counting <= '0'5��    <   "                  G                     5�_�   �   �           �   >   #    ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f�     �   =   ?   �      #            elsif is_counting = '1'5��    =   #                  l                     �    =   )                  r                     �    =   (                  q                     �    =   '                 p                    �    =   '                 p                    �    =   '                 p                    �    =   +                  t                     �    =   *                  s                     �    =   )                  r                     �    =   (                  q                     �    =   '                  p                     5�_�   �   �           �   >   '    ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f�      �   =   ?   �      '            elsif is_counting = '1' or 5��    =   '                  p                     5�_�   �   �           �   >   (    ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f�      �   =   ?   �      )            elsif is_counting = '1' or ()5��    =   (                  q                     �    =   (                 q                    �    =   (                 q                    �    =   (                 q                    5�_�   �   �           �   >   0    ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f�#     �   =   ?   �      1            elsif is_counting = '1' or (start = )5��    =   0                  y                     5�_�   �   �           �   >   1    ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f�$     �   =   ?   �      3            elsif is_counting = '1' or (start = '')5��    =   1                  z                     �    =   1                 z                    5�_�   �   �           �   >   3    ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f�&     �   =   ?   �      4            elsif is_counting = '1' or (start = '0')5��    =   3               	   |              	       �    =   8                 �                    �    =   8                 �                    �    =   8                 �                    �    =   8                 �                    �    =   8              
   �             
       5�_�   �   �           �   >   B    ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f�4     �   =   ?   �      C            elsif is_counting = '1' or (start = '0' and counter = )5��    =   B                  �                     5�_�   �   �           �   >   C    ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f�4     �   =   ?   �      E            elsif is_counting = '1' or (start = '0' and counter = '')5��    =   C                  �                     5�_�   �   �           �   >   F    ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f�6     �   =   ?   �      F            elsif is_counting = '1' or (start = '0' and counter = '0')5��    =   F                  �                     5�_�   �   �           �   >   C    ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f�y     �   =   ?   �      K            elsif is_counting = '1' or (start = '0' and counter = '0') then5��    =   C                 �                    5�_�   �   �           �   >   C    ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f�{     �   =   ?   �      K            elsif is_counting = '1' or (start = '0' and counter = '1') then5��    =   C                 �                    5�_�   �   �           �   >   8    ����                                                                                                                                                                                                                                                                                                                            ~          |          V       f�     �   =   ?   �      K            elsif is_counting = '1' or (start = '0' and counter = '0') then5��    =   8                 �                    �    =   9                  �                     �    =   8                 �                    �    =   8                 �                    �    =   8                 �                    5�_�   �   �           �   ?   &    ����                                                                                                                                                                                                                                                                                                                            ~          |          V       fы     �   ?   A   �                      �   ?   A   �    5��    ?                      �                     �    ?                     �                     �    ?                     �                     �    ?                    �                    �    ?                    �                    �    ?                    �                    �    ?                    �                    5�_�   �   �           �   @       ����                                                                                                                                                                                                                                                                                                                                      }          V       fё     �   ?   A   �                      is_counting <= 5��    ?                     �                     5�_�   �   �           �   @        ����                                                                                                                                                                                                                                                                                                                                      }          V       fђ     �   ?   A   �      !                is_counting <= ''5��    ?                      �                     5�_�   �   �           �   @   "    ����                                                                                                                                                                                                                                                                                                                                      }          V       fѓ    �   ?   A   �      "                is_counting <= '1'5��    ?   "                  �                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�u     �   �   �       S   (architecture Behavioral of serial_out is       type state_t is (           INICIO, START_BIT,   i        TRANSMISSAO0, TRANSMISSAO1, TRANSMISSAO2, TRANSMISSAO3, TRANSMISSAO4, TRANSMISSAO5, TRANSMISSAO6,           STOP_BIT   
        );   +    signal estado_atual: state_t := INICIO;   ,    signal prox_estado: state_t:= START_BIT;   "    signal enviados: integer := 0;           p1: process(clk) begin   "        if (rising_edge(clk)) then   (            estado_atual <= prox_estado;           end if;               if (reset = '1') then   #            estado_atual <= INICIO;   "            prox_estado <= INICIO;               enviados <= 0;           end if;               case estado_atual is                when INICIO =>                   tx_done <= '0';                    serial_o <= '1';                   enviados <= 0;   #                if tx_go = '1' then   -                    prox_estado <= START_BIT;                   else       *                    prox_estado <= INICIO;                   end if;                   when START_BIT =>                   tx_done <= '0';                    serial_o <= '0';   ,                prox_estado <= TRANSMISSAO0;                               when TRANSMISSAO0 =>                   tx_done <= '0';   $                serial_o <= data(0);   ,                prox_estado <= TRANSMISSAO1;                               when TRANSMISSAO1 =>                   tx_done <= '0';   $                serial_o <= data(1);   ,                prox_estado <= TRANSMISSAO2;                               when TRANSMISSAO2 =>                   tx_done <= '0';   $                serial_o <= data(2);   ,                prox_estado <= TRANSMISSAO3;                               when TRANSMISSAO3 =>                   tx_done <= '0';   $                serial_o <= data(3);   ,                prox_estado <= TRANSMISSAO4;                    when TRANSMISSAO4 =>                   tx_done <= '0';   $                serial_o <= data(4);   ,                prox_estado <= TRANSMISSAO5;                    when TRANSMISSAO5 =>                   tx_done <= '0';   $                serial_o <= data(5);   ,                prox_estado <= TRANSMISSAO6;                    when TRANSMISSAO6 =>                   tx_done <= '0';   $                serial_o <= data(6);   (                prox_estado <= STOP_BIT;                              when STOP_BIT =>                   tx_done <= '1';                    serial_o <= '1';   &                prox_estado <= INICIO;                   when others =>   &                prox_estado <= INICIO;               end case;       end process p1;   end architecture;    5��    �       S               �      �	              5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        f�~     �   �   �   �      !    done <= '1' when reset = '1';       lg: process(clock, reset)   	    begin           if reset = '1' then               done <= '1';               tx_done <= '1';               is_counting <= '0';   %        elsif rising_edge(clock) then   /            if i = 0 and is_counting = '0' then               end if;       end process lg;5��    �                     �      6      ]      5�_�   �   �           �   {        ����                                                                                                                                                                                                                                                                                                                            �           �           V        fӁ     �   z   |   �      3        port map(clock, reset, not is_counting, i);5��    z                           4       7       5�_�   �   �           �   y        ����                                                                                                                                                                                                                                                                                                                            z           y           V        fӅ    �   x   {   �      !    data_counter: counter_generic   a        generic map(WIDTH+2+STOP_BITS)    -- The sums are to send the start, parity and stop bits5��    x                     �
      �       �       5�_�   �   �   �       �   /       ����                                                                                                                                                                                                                                                                                                                            z           y           V        f��     �   .   0   �          signal counter: natural;5��    .                     �                     5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            z           y           V        f��     �   /   1   �          signal is_counting: bit;5��    /                                          5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            z           y           V        f��     �   /   1   �           signal is_counting: bit := ;5��    /                                          5�_�   �   �           �   0        ����                                                                                                                                                                                                                                                                                                                            z           y           V        f��   	 �   /   1   �      "    signal is_counting: bit := '';5��    /                                           5�_�   �   �           �   :        ����                                                                                                                                                                                                                                                                                                                            z           y           V        f�Z     �   :   <   �                  �   :   <   �    5��    :                      �              	       �    :                     �                    5�_�   �   �           �   ;       ����                                                                                                                                                                                                                                                                                                                            {           z           V        f�_     �   :   <   �                  report 5��    :                     �                     5�_�   �   �           �   ;       ����                                                                                                                                                                                                                                                                                                                            {           z           V        f�a     �   :   <   �                  report ""5��    :                     �                     5�_�   �   �           �   ;       ����                                                                                                                                                                                                                                                                                                                            {           z           V        f�d     �   :   <   �                  report "";5��    :                     �                     �    :                 
                
       5�_�   �   �           �   ;   #    ����                                                                                                                                                                                                                                                                                                                            {           z           V        f�n     �   :   <   �      $            report "counter is in ";5��    :   #                                       5�_�   �   �           �   ;   3    ����                                                                                                                                                                                                                                                                                                                            {           z           V        f�w     �   :   <   �      4            report "counter is in " & integer'image;5��    :   3                                       5�_�   �   �           �   ;   4    ����                                                                                                                                                                                                                                                                                                                            {           z           V        f�x   
 �   :   <   �      6            report "counter is in " & integer'image();5��    :   4                                       �    :   8                 "                    5�_�   �   �   �       �   ;       ����                                                                                                                                                                                                                                                                                                                            {           z           V        f՝    �   :   <   �      =            report "counter is in " & integer'image(counter);5��    :                     �                     5�_�   �   �           �   ;       ����                                                                                                                                                                                                                                                                                                                            {           z           V        fխ     �   :   ;          J            assert false report "counter is in " & integer'image(counter);5��    :                      �      K               5�_�   �   �   �       �   >       ����                                                                                                                                                                                                                                                                                                                            >          >   I       v   I    f�`     �   =   ?   �      O            elsif is_counting = '1' or (start = '0' and is_counting = '0') then5��    =                     a                     5�_�   �   �           �   >       ����                                                                                                                                                                                                                                                                                                                            >          >   I       v   I    f�`     �   =   ?   �      N            lsif is_counting = '1' or (start = '0' and is_counting = '0') then5��    =                     a                     5�_�   �   �           �   >       ����                                                                                                                                                                                                                                                                                                                            >          >   I       v   I    f�a     �   =   ?   �      M            sif is_counting = '1' or (start = '0' and is_counting = '0') then5��    =                     a                     5�_�   �   �           �   >       ����                                                                                                                                                                                                                                                                                                                            >          >   I       v   I    f�d    �   =   ?   �    �   >   ?   �    5��    =                      U                     5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                                                             f�I     �   -   /   �      &architecture rtl of counter_generic is5��    -                    �                    �    -                    �                    �    -                    �                    �    -                 
   �             
       �    -          
       
   �      
       
       �    -          
          �      
              �    -                 
   �             
       5�_�   �   �           �   H       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   G   I   �      end architecture rtl;5��    G                     s                     5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                                                             f�S     �   .   0   �      !    signal counter: natural := 0;5��    .                                        �    .                                        �    .                                           �    .                 	                	       �    .          	                	              �    .                                        5�_�   �   �           �   7       ����                                                                                                                                                                                                                                                                                                                                                             f�i     �   6   8   �                  counter <= 0;5��    6                    �                    �    6                     �                     �    6                    �                    �    6                     �                     �    6                     �                     �    6                 	   �             	       �    6          	          �      	              �    6                    �                    �    6                    �                    �    6                    �                    5�_�   �   �           �   8       ����                                                                                                                                                                                                                                                                                                                                                             f�4     �   7   9   �                  done <= '0';5��    7                     �                     �    7                     �                     �    7                     �                     5�_�   �   �           �   8       ����                                                                                                                                                                                                                                                                                                                                                             f�7     �   7   9   �                  done <= ;5��    7                     �                     5�_�   �   �           �   8       ����                                                                                                                                                                                                                                                                                                                                                             f�9     �   7   9   �                  done <= '';5��    7                     �                     5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                                                             f�Q     �   /   0          #    signal is_counting: bit := '0';5��    /                            $               5�_�   �   �           �   8        ����                                                                                                                                                                                                                                                                                                                                                             f�V     �   7   8                      is_counting <= '0';5��    7                      �                      5�_�   �   �           �   ;        ����                                                                                                                                                                                                                                                                                                                                                             f�X     �   :   ;          #                is_counting <= '0';5��    :                            $               5�_�   �   �           �   >       ����                                                                                                                                                                                                                                                                                                                                                             f�]     �   =   >          #                is_counting <= '1';5��    =                      �      $               5�_�   �   �           �   <       ����                                                                                                                                                                                                                                                                                                                            <          <   F       v   F    f�q     �   ;   =   �      L            if is_counting = '1' or (start = '0' and is_counting = '0') then5��    ;          8          +      8              �    ;                     -                     �    ;                     ,                     �    ;                    +                    �    ;                     .                     �    ;                     -                     �    ;                     ,                     �    ;                    +                    �    ;                    +                    �    ;                    +                    �    ;                     6                     �    ;                    5                    �    ;                    5                    �    ;                    5                    5�_�   �   �           �   <       ����                                                                                                                                                                                                                                                                                                                            <          <   F       v   F    f��     �   ;   =   �      )            if counter < MAX_COUNT-1 then5��    ;                     +                     5�_�   �   �           �   <       ����                                                                                                                                                                                                                                                                                                                            <          <   F       v   F    f��     �   ;   =   �      *            if (counter < MAX_COUNT-1 then5��    ;                           +       ,       5�_�   �              �   <   &    ����                                                                                                                                                                                                                                                                                                                            <          <   F       v   F    f��     �   ;   =   �      +            if (counter < MAX_COUNT-1) then5��    ;   &                  B                     5�_�   �                <   *    ����                                                                                                                                                                                                                                                                                                                            <          <   F       v   F    f��     �   ;   =   �      /            if (counter < MAX_COUNT-1) or  then5��    ;   *                  F                     5�_�                  <   +    ����                                                                                                                                                                                                                                                                                                                            <          <   F       v   F    f��     �   ;   =   �      1            if (counter < MAX_COUNT-1) or () then5��    ;   +                  G                     �    ;   +                 G                    �    ;   +                 G                    �    ;   +                 G                    5�_�                 <   3    ����                                                                                                                                                                                                                                                                                                                            <          <   F       v   F    f��     �   ;   =   �      9            if (counter < MAX_COUNT-1) or (start = ) then5��    ;   3                  O                     5�_�                 <   4    ����                                                                                                                                                                                                                                                                                                                            <          <   F       v   F    f��     �   ;   =   �      ;            if (counter < MAX_COUNT-1) or (start = '') then5��    ;   4                  P                     5�_�                 <   6    ����                                                                                                                                                                                                                                                                                                                            <          <   F       v   F    f��    �   ;   =   �      <            if (counter < MAX_COUNT-1) or (start = '1') then5��    ;   6               	   R              	       �    ;   >                  Z                     �    ;   =                  Y                     �    ;   <                  X                     �    ;   ;                 W                    �    ;   ;                 W                    �    ;   ;                 W                    �    ;   E                 a                    �    ;   F                  b                     �    ;   E                 a                    �    ;   G                  c                     �    ;   F                  b                     �    ;   E                 a                    �    ;   E                 a                    �    ;   E                 a                    �    ;   E                 a                    5�_�                 6       ����                                                                                                                                                                                                                                                                                                                            9   (       9   (       V   O    f��     �   5   7   �      #            counter <= MAX_COUNT-1;5��    5                    w                    5�_�                 :       ����                                                                                                                                                                                                                                                                                                                            9   (       9   (       V   O    f��     �   :   <   �                      �   :   <   �    5��    :                      �                     �    :                                          �    :                                          �    :                                          �    :                                        �    :                                        �    :                                        5�_�                 =       ����                                                                                                                                                                                                                                                                                                                            9   (       9   (       V   O    f�     �   <   >   �      V            if (counter < MAX_COUNT-1) or (start = '1' and counter = MAX_COUNT-1) then5��    <                    H                    5�_�    	             =       ����                                                                                                                                                                                                                                                                                                                            9   (       9   (       V   O    f�     �   <   >   �      V            if (counter > MAX_COUNT-1) or (start = '1' and counter = MAX_COUNT-1) then5��    <                    J                    5�_�    
          	   =       ����                                                                                                                                                                                                                                                                                                                            9   (       9   (       V   O    f�)     �   <   >   �      L            if (counter > 0) or (start = '1' and counter = MAX_COUNT-1) then5��    <                     K                     �    <   !                  Q                     �    <                      P                     �    <                     O                     �    <                     N                     �    <                     M                     �    <                     K                     5�_�  	            
   =   ;    ����                                                                                                                                                                                                                                                                                                                            9   (       9   (       V   O    f�A    �   <   >   �      L            if (counter > 0) or (start = '1' and counter = MAX_COUNT-1) then5��    <   ;                 k                    5�_�  
               /       ����                                                                                                                                                                                                                                                                                                                                        E           V        f    �   .   0   �      +    signal counter: natural := MAX_COUNT-1;5��    .                                        5�_�                 3       ����                                                                                                                                                                                                                                                                                                                                        E           V        f&�    �   2   4   �          counting: process(clk, rst)5��    2                     0                     �    2   "                  4                     �    2   !                  3                     �    2                     2                    �    2                     2                    �    2                     2                    5�_�                          ����                                                                                                                                                                                                                                                                                                                                        E           V        f�l    �              &   library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity counter_generic is       generic(           MAX_COUNT: natural       );   
    port (   J        clk, rst, start: in bit;                            -- Clock input           done: out bit;   B        count : out natural       -- 6-bit count output (64 steps)       );   end counter_generic;       -architecture Behavioral of counter_generic is   !    signal counter: natural := 0;       begin          &    counting: process(clk, rst, start)   	    begin           if rst = '1' then               counter <= 0;               done <= '0';   #        elsif rising_edge(clk) then   )            if counter = MAX_COUNT-1 then                   done <= '1';                   counter <= 0;               end if;   B            if (counter > 0) or (start = '1' and counter = 0) then   '                counter <= counter + 1;               end if;           end if;       end process counting;           count <= counter;          end architecture;5��           &               w      �              5�_�                 4       ����                                                                                                                                                                                                                                                                                                                                                             fĨ     �   3   5   g      (architecture Behavioral of serial_out is5��    3          
                
              5�_�                 f       ����                                                                                                                                                                                                                                                                                                                                                             fĮ     �   e   g   g      end architecture Behavioral;5��    e          
           <	      
               5�_�                 f       ����                                                                                                                                                                                                                                                                                                                                                             fĮ    �   e   g   g      end architecture ;5��    e                     ;	                     5�_�                 %       ����                                                                                                                                                                                                                                                                                                                                                             fƿ     �   $   &   g      entity serial_out is5��    $                     �                     5�_�                 2       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   1   3   g      end serial_out;5��    1                                          5�_�                 4       ����                                                                                                                                                                                                                                                                                                                                                             f��     �   3   5   g      !architecture rtl of serial_out is5��    3                     0                     5�_�                 4        ����                                                                                                                                                                                                                                                                                                                                                             f��     �   3   5   g      $architecture rtl of serial_out_v) is5��    3                     2                    5�_�                 4        ����                                                                                                                                                                                                                                                                                                                                                             f��    �   3   5   g      $architecture rtl of serial_out_v) is5��    3                     2                    5�_�                          ����                                                                                                                                                                                                                                                                                                                            g                     V   /    f�
    �               g   library IEEE;   use IEEE.NUMERIC_BIT.all;       entity generic_reg is       generic(           WIDTH: natural := 8       );   
    port (   !        rst, clk, enable: in bit;   +        d: in bit_vector(WIDTH-1 downto 0);   +        q: out bit_vector(WIDTH-1 downto 0)       );   end entity generic_reg;       'architecture Behavior of generic_reg is   /    signal value: bit_vector(WIDTH-1 downto 0);   begin              process(rst, clk)   	    begin           if rst = '1' then   %            value <= (others => '0');   4        elsif rising_edge(clk) and enable = '1' then               value <= D;           end if;       end process;           q <= value;          end architecture Behavior;           -- 8 bits de dados   library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity serial_out_V0 is       generic(   #        POLARITY : boolean := TRUE;           WIDTH: natural := 7;           PARITY : natural := 1;            STOP_BITS : natural := 1       );   	    port(   %        clock, reset, tx_go : in bit;           tx_done : out bit;   /        data : in bit_vector(WIDTH-1 downto 0);           serial_o : out bit       );   end serial_out_v0;       $architecture rtl of serial_out_v0 is           component generic_reg           generic(               WIDTH: natural   
        );           port (   %            rst, clk, enable: in bit;   /            d: in bit_vector(WIDTH-1 downto 0);   /            q: out bit_vector(WIDTH-1 downto 0)   
        );       end component;           component counter_generic           generic(               MAX_COUNT: natural   
        );           port (   N            clk, rst, start: in bit;                            -- clock input               done: out bit;   F            count : out natural       -- 6-bit count output (64 steps)   
        );       end component;           signal i: natural;       signal done: bit;          begin       $    -- data_counter: counter_generic   d    --     generic map(WIDTH+2+STOP_BITS)    -- The sums are to send the start, parity and stop bits   6        -- port map(clock, reset, not is_counting, i);       "    -- counting_state: generic_reg       --     generic map(1)   #    --     port map(reset, clock, )       $    -- done <= '1' when reset = '1';        -- lg: process(clock, reset)       -- begin       --     if reset = '1' then       --         done <= '1';       --         tx_done <= '1';   "    --         is_counting <= '0';   (    --     elsif rising_edge(clock) then   2    --         if i = 0 and is_counting = '0' then       --       --     end if;       -- end process lg;          end architecture;    5��            g       g               G	      n
      5�_�   �           �   �   >       ����                                                                                                                                                                                                                                                                                                                            >          >   I       v   I    f�8     �   =   ?   �                  elsif  then5��    =          8           g      8               5�_�   �           �   �   ;   :    ����                                                                                                                                                                                                                                                                                                                            z           y           V        fՎ     �   :   <        5��    :                      �      >               5�_�   �   �       �   �      .    ����                                                                                                                                                                                                                                                                                                                            z           y           V        f��     �         �      3    signal value: bit_vector(WIDTH-1 downto 0) := ;5��       .                  j                     5�_�   �   �           �      2    ����                                                                                                                                                                                                                                                                                                                            z           y           V        f��     �         �      5    signal value: bit_vector(WIDTH-1 downto 0) := ();5��       2                  n                     5�_�   �               �      3    ����                                                                                                                                                                                                                                                                                                                            z           y           V        f��     �         �      B    signal value: bit_vector(WIDTH-1 downto 0) := (others => '0');5��       3                  o                     �       3                 o                    �       3                 o                    �       3                 o                    �       3                 o                    5�_�   �           �   �   u       ����                                                                                                                                                                                                                                                                                                                            |          |          v       f2�     �   t   u   �       5��    t                      �	                     �    t                      �	                     5�_�   Z           \   [   P       ����                                                                                                                                                                                                                                                                                                                            9          9   !       v       f,�     �   O   Q   �      
    port (5��    O                     y                     5�_�   K           M   L   [        ����                                                                                                                                                                                                                                                                                                                            [          [                 f+�     �   Z   f        5��    Z                      G                    5�_�   0           2   1   3   %    ����                                                                                                                                                                                                                                                                                                                            3          3   &       v       f�     �   2   4   �      7            if to_integer(counter) = others => '0' then5��    2   %                 �                    �    2   %                 �                    �    2   %                 �                    �    2   %                 �                    �    2   %                 �                    5�_�   +           -   ,   5       ����                                                                                                                                                                                                                                                                                                                            4          4   &       v       fo     �   4   5   �                      �   4   6   �                      don5��    4                      �                     �    4                     �                    5�_�                     3       ����                                                                                                                                                                                                                                                                                                                            2          2          v   %    fD     �   3   4   �    �   2   4   �      0            donto_integer(counter) = 63e <= '1';5��    2                     y                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       fG     �      	   �      $       d: in bit_vector(7 downto 0);5��                          �                      5��