Vim�UnDo� ��~T}@u���/@���Ǹղ�U���Ȳ�   G   6            " X=" & 'image(to_integer(signed(x))) &LF&   8                    e��   9 _�                             ����                                                                                                                                                                                                                                                                                                                                                             e�L�     �                   �               5��                                                  �                                                �                                                �                                                  �                    H                       R      5�_�                            ����                                                                                                                                                                                                                                                                                                                                       I           V        e�Mq     �                  library IEEE;�               �             H   use IEEE.STD_LOGIC_1164.ALL;   use IEEE.STD_LOGIC_ARITH.ALL;    use IEEE.STD_LOGIC_UNSIGNED.ALL;       entity ch_test is   end entity ch_test;       $architecture testbench of ch_test is       -- Constants   (    constant CLK_PERIOD : time := 10 ns;            -- Signals for the testbench   6    signal x_tb, y_tb, z_tb : bit_vector(31 downto 0);   @    signal q_tb_expected, q_tb_actual : bit_vector(31 downto 0);       <    -- Component declaration for the DUT (Design Under Test)       component ch           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;       begin       -- Instantiate the DUT       DUT_inst : ch   E        port map (x => x_tb, y => y_tb, z => z_tb, q => q_tb_actual);           -- Stimulus process       stimulus_process: process   	    begin           -- Test case 1            x_tb <= (others => '0');            y_tb <= (others => '1');            z_tb <= (others => '0');           wait for CLK_PERIOD;                      -- Test case 2            x_tb <= (others => '1');            y_tb <= (others => '0');            z_tb <= (others => '1');           wait for CLK_PERIOD;       (        -- Add more test cases as needed       A        wait; -- Wait indefinitely to keep the simulation running       end process;           -- Check results process   "    check_results_process: process   	    begin   L        wait for 2 * CLK_PERIOD; -- Allow time for the DUT to produce output                      -- Test case 1   )        q_tb_expected <= (others => '0');   *        assert q_tb_actual = q_tb_expected   '            report "Test case 1 failed"               severity failure;               -- Test case 2   )        q_tb_expected <= (others => '1');   *        assert q_tb_actual = q_tb_expected   '            report "Test case 2 failed"               severity failure;       G        -- Add more result checking as needed for additional test cases               wait;       end process;       end testbench;    5��           H                      E              �                                                  �                    A                       $      5�_�                            ����                                                                                                                                                                                                                                                                                                                                       B           V        e�N
     �                  library IEEE;�               �             A   use IEEE.STD_LOGIC_1164.ALL;   use IEEE.STD_LOGIC_ARITH.ALL;    use IEEE.STD_LOGIC_UNSIGNED.ALL;       entity ch_test is   end entity ch_test;       $architecture testbench of ch_test is       -- Constants   (    constant CLK_PERIOD : time := 10 ns;            -- Type for test case vector   !    type test_case_type is record   <        x_value, y_value, z_value : bit_vector(31 downto 0);   -        q_expected : bit_vector(31 downto 0);       end record;           -- Vector of test cases   <    constant test_cases : array(0 to 1) of test_case_type :=   	        (   �            (x_value => (others => '0'), y_value => (others => '1'), z_value => (others => '0'), q_expected => (others => '0')),               (x_value => (others => '1'), y_value => (others => '0'), z_value => (others => '1'), q_expected => (others => '1'))   ,            -- Add more test cases as needed   
        );            -- Signals for the testbench   6    signal x_tb, y_tb, z_tb : bit_vector(31 downto 0);   @    signal q_tb_expected, q_tb_actual : bit_vector(31 downto 0);       <    -- Component declaration for the DUT (Design Under Test)       component ch           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;       begin       -- Instantiate the DUT       DUT_inst : ch   E        port map (x => x_tb, y => y_tb, z => z_tb, q => q_tb_actual);           -- Testbench process       testbench_process: process   	    begin   &        for i in test_cases'range loop   9            -- Set input values for the current test case   *            x_tb <= test_cases(i).x_value;   *            y_tb <= test_cases(i).y_value;   *            z_tb <= test_cases(i).z_value;       L            wait for CLK_PERIOD; -- Allow time for the DUT to produce output       5            -- Check result for the current test case   6            q_tb_expected <= test_cases(i).q_expected;   .            assert q_tb_actual = q_tb_expected   B                report "Test case " & integer'image(i) & " failed"   !                severity failure;           end loop;       A        wait; -- Wait indefinitely to keep the simulation running       end process;       end testbench;    5��           A                                    �                                                  �                    H                             5�_�                            ����                                                                                                                                                                                                                                                                                                                                       J           V        e�N    �                  library IEEE;�               �             H   use IEEE.STD_LOGIC_1164.ALL;   use IEEE.STD_LOGIC_ARITH.ALL;    use IEEE.STD_LOGIC_UNSIGNED.ALL;       entity ch_test is   end entity ch_test;       $architecture testbench of ch_test is       -- Constants   (    constant CLK_PERIOD : time := 10 ns;            -- Signals for the testbench   6    signal x_tb, y_tb, z_tb : bit_vector(31 downto 0);   @    signal q_tb_expected, q_tb_actual : bit_vector(31 downto 0);       <    -- Component declaration for the DUT (Design Under Test)       component ch           port (   0            x, y, z: in bit_vector(31 downto 0);   *            q: out bit_vector(31 downto 0)   
        );       end component;           -- Vector of test cases   Q    type test_vector_type is array (natural range <>) of bit_vector(31 downto 0);   0    constant test_vector : test_vector_type := (   (        (others => '0'),  -- Test case 1   (        (others => '1')   -- Test case 2   (        -- Add more test cases as needed       );       begin       -- Stimulus process       stimulus_process: process   	    begin   '        for i in test_vector'range loop   ?            -- Apply the input vector for the current test case   #            x_tb <= test_vector(i);   $            y_tb <= (others => '1');   $            z_tb <= (others => '0');                               wait for CLK_PERIOD;       C            -- Add more stimuli as needed for the current test case           end loop;       A        wait; -- Wait indefinitely to keep the simulation running       end process;           -- Check results process   "    check_results_process: process   	    begin   '        for i in test_vector'range loop   7            -- Allow time for the DUT to produce output                wait for CLK_PERIOD;       B            -- Apply the expected output for the current test case   -            q_tb_expected <= (others => '0');   .            assert q_tb_actual = q_tb_expected   F                report "Test case " & integer'image(i + 1) & " failed"   !                severity failure;       K            -- Add more result checking as needed for the current test case           end loop;               wait;       end process;           -- Instantiate the DUT       DUT_inst : ch           port map (x => x_    5��           H                                    �                                                  �                    J                       T      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       e�PJ    �                use IEEE.STD_LOGIC_1164.ALL;   use IEEE.STD_LOGIC_ARITH.ALL;    use IEEE.STD_LOGIC_UNSIGNED.ALL;5��                                 \               5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       e�P�     �         G              �         G    �         G      0    constant test_vector : test_vector_type := (    �         G      (        (others => '0'),  -- Test case 1�                (        (others => '1')   -- Test case 25��                          �      )               �                          �                      �                         �                    �                          �                     �                          �                     �                          �                     �                          �                     �                          �                     �       0                  �                     �       0                 �                     �                         �                     �                     <   �              ,      5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                       e�Q     �         K      <    (x"00000001", x"00000002", x"00000004"),  -- Test case 3   <    (x"AAAA5555", x"5555AAAA", x"AAAA5555"),  -- Test case 4   <    (x"12345678", x"87654321", x"13579BDF"),  -- Test case 5�         K      <    (x"FFFFFFFF", x"00000000", x"FFFFFFFF"),  -- Test case 25��                         �                     �                         -                     �                         n                     �                         �                     5�_�      
          	      /    ����                                                                                                                                                                                                                                                                                                                                                       e�Q    �         K      @        (x"12345678", x"87654321", x"13579BDF"),  -- Test case 55��       /                  �                     5�_�   	              
   '       ����                                                                                                                                                                                                                                                                                                                            '   !       '          v       e�Q9     �   &   (   K      #            x_tb <= test_vector(i);�   '   (   K    5��    &                    �                    5�_�   
                 (       ����                                                                                                                                                                                                                                                                                                                            (          )   "          "    e�QE    �   '   )   K                  y_tb <= ;�   (   )   K    �   '   *   K      $            y_tb <= (others => '1');   $            z_tb <= (others => '0');5��    '                                          �    (                     %                     �    '                                          �    (                     @                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            (          (   .          "    e��     �         K      end entity ch_test;5��                         %                      5�_�                           ����                                                                                                                                                                                                                                                                                                                            (          (   .          "    e��     �         K      end ;5��                         $                      5�_�                            ����                                                                                                                                                                                                                                                                                                                            (          (   .          "    e��    �         K      entity ch_test is   end;�         K      end;5��                                                �                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                            '          '   .          "    e�     �         J      $architecture testbench of ch_test is5��              	          4       	              5�_�                    I       ����                                                                                                                                                                                                                                                                                                                            '          '   .          "    e�     �   H   J   J      end testbench;5��    H          	          �      	              �    H                     �                     �    H                    �                    �    H                    �                    �    H                    �                    5�_�                    E        ����                                                                                                                                                                                                                                                                                                                            E          H           V       e�     �   D   E              -- Instantiate the DUT       DUT_inst : ch   E        port map (x => x_tb, y => y_tb, z => z_tb, q => q_tb_actual);    5��    D                      w      t               5�_�                            ����                                                                                                                                                                                                                                                                                                                            E          E           V       e�*     �       %   F    �       !   F    5��                                         t       5�_�                    &       ����                                                                                                                                                                                                                                                                                                                            I          I           V       e     �   %   '   J          stimulus_process: process5��    %                     �                     �    %                     �                    5�_�                    &       ����                                                                                                                                                                                                                                                                                                                            I          I           V       e     �   %   '   J      .                  stimulus_process: process is5��    %                     �                     5�_�                    &       ����                                                                                                                                                                                                                                                                                                                            I          I           V       e     �   %   '   J           stimulus_process: process is5��    %                    �                    5�_�                            ����                                                                                                                                                                                                                                                                                                                            I          I           V       e�P/     �          J      library IEEE;�         J    5��                                                  �                                           "       5�_�                            ����                                                                                                                                                                                                                                                                                                                            K          K           V       e�P0     �                 5��                          "                      5�_�                   '       ����                                                                                                                                                                                                                                                                                                                            J          J           V       e�Pe     �   '   -   L              �   (   )   L    �   '   )   K    5��    '                      �                     �    '                     �                    �    '                     �              �       5�_�                    '       ����                                                                                                                                                                                                                                                                                                                            O          O           V       e�Ph     �   &   (   P          st: process is5��    &                    �                    5�_�                    (   
    ����                                                                                                                                                                                                                                                                                                                            O          O           V       e�Pk     �   '   )   P      =          file tb_file : text open read_mode is "alu_tb.dat";5��    '                     �                     5�_�                    )       ����                                                                                                                                                                                                                                                                                                                            )          +                 e�Po    �   )   ,   P        variable space: character;   0  variable Av, Bv, res: bit_vector(63 downto 0);�   (   *   P        variable tb_line: line;5��    (                                           �    )                                           �    *                     C                     5�_�                    (   /    ����                                                                                                                                                                                                                                                                                                                            )          +                 e�P�   	 �   '   )   P      ;        file tb_file : text open read_mode is "alu_tb.dat";5��    '   /       
       	   �      
       	       5�_�                     +       ����                                                                                                                                                                                                                                                                                                                            )          +                 e�P�     �   *   ,   P      6        variable Av, Bv, res: bit_vector(63 downto 0);5��    *                    Q                    �    *                    Q                    �    *                    Q                    �    *                    Q                    5�_�      !               +       ����                                                                                                                                                                                                                                                                                                                            )          +                 e�P�     �   *   ,   P      8        variable x_tb, Bv, res: bit_vector(63 downto 0);5��    *                    W                    �    *                    W                    �    *                    W                    �    *                    W                    5�_�       "           !   +       ����                                                                                                                                                                                                                                                                                                                            )          +                 e�P�     �   *   ,   P      :        variable x_tb, y_tb, res: bit_vector(63 downto 0);5��    *                     \                     �    *                    ]                    �    *                    ]                    �    *                    ]                    5�_�   !   #           "   +   3    ����                                                                                                                                                                                                                                                                                                                            )          +                 e�P�   
 �   *   ,   P      @        variable x_tb, y_tb, z_tb, res: bit_vector(63 downto 0);5��    *   3                 s                    5�_�   "   %           #   /        ����                                                                                                                                                                                                                                                                                                                            .   &       7          V   4    e�S!     �   -   7   G      '        for i in test_vector'range loop�   .   /   G    �   .   /       	   ?            -- Apply the input vector for the current test case   0            x_tb <= test_vector(i)(31 downto 0);   0            y_tb <= test_vector(i)(31 downto 0);   0            z_tb <= test_vector(i)(31 downto 0);                               wait for CLK_PERIOD;       C            -- Add more stimuli as needed for the current test case           end loop;5��    .       	               �      X              �    -                     �                     �    -                     �              �       5�_�   #   &   $       %   /       ����                                                                                                                                                                                                                                                                                                                            /          5                 e�SA     �   /   6   O        readline(tb_file, tb_line);     read(tb_line, Av);     A <= signed(Av);     read(tb_line, space);     read(tb_line, Bv);     B <= signed(Bv);�   .   0   O        -- read inputs5��    .                  
   �              
       �    /                  
   �              
       �    0                  
   �              
       �    1                  
                 
       �    2                  
   5              
       �    3                  
   W              
       �    4                  
   v              
       5�_�   %   '           &   +        ����                                                                                                                                                                                                                                                                                                                            +          +          V       e�S^     �   *   ,   O      @        variable x_tb, y_tb, z_tb, res: bit_vector(31 downto 0);5��    *                    S                    �    *                    X                    �    *                    ]                    5�_�   &   (           '   +       ����                                                                                                                                                                                                                                                                                                                            +          +          V       e�S     �   *   ,   O      =        variable x_v, y_v, z_v, res: bit_vector(31 downto 0);5��    *                    Q                    5�_�   '   )           (   +       ����                                                                                                                                                                                                                                                                                                                            +          +          V       e�S�     �   *   ,   O      <        variable Xv, y_v, z_v, res: bit_vector(31 downto 0);5��    *                    U                    5�_�   (   *           )   +       ����                                                                                                                                                                                                                                                                                                                            +          +          V       e�S�     �   *   ,   O      ;        variable Xv, Yv, z_v, res: bit_vector(31 downto 0);5��    *                    Y                    5�_�   )   +           *   1       ����                                                                                                                                                                                                                                                                                                                            +          +          V       e�S�     �   0   2   O                  read(tb_line, Av);5��    0                                        5�_�   *   ,           +   2       ����                                                                                                                                                                                                                                                                                                                            +          +          V       e�S�     �   1   3   O                  A <= signed(Av);5��    1                    (                    5�_�   +   -           ,   2       ����                                                                                                                                                                                                                                                                                                                            +          +          V       e�S�     �   1   3   O                  A <= signed(Xv);5��    1                                        5�_�   ,   .           -          ����                                                                                                                                                                                                                                                                                                                            +          +          V       e��v     �         O      entity ch_test is end;5��                        .                     5�_�   -   /           .          ����                                                                                                                                                                                                                                                                                                                            +          +          V       e��|     �         O      architecture dut of ch_test is5��                        Q                     5�_�   .   0           /   #       ����                                                                                                                                                                                                                                                                                                                            +          +          V       e���     �   "   $   O          DUT_inst : ch5��    "                    <                    5�_�   /   1           0   #       ����                                                                                                                                                                                                                                                                                                                            +          +          V       e���     �   "   $   O          dut : ch5��    "                     ?                     5�_�   0   2           1           ����                                                                                                                                                                                                                                                                                                                                                  V       e���     �                    -- Vector of test cases   Q    type test_vector_type is array (natural range <>) of bit_vector(31 downto 0);   0    constant test_vector : test_vector_type := (   @        (x"00000000", x"00000000", x"00000000"),  -- Test case 1   @        (x"FFFFFFFF", x"00000000", x"FFFFFFFF"),  -- Test case 2   @        (x"00000001", x"00000002", x"00000004"),  -- Test case 3   @        (x"AAAA5555", x"5555AAAA", x"AAAA5555"),  -- Test case 4   ?        (x"12345678", x"87654321", x"13579BDF")  -- Test case 5   (        -- Add more test cases as needed       );    5��                                              5�_�   1   3           2           ����                                                                                                                                                                                                                                                                                                                                                V       e��F     �                @    signal q_tb_expected, q_tb_actual : bit_vector(31 downto 0);�   
      D      6    signal x_tb, y_tb, z_tb : bit_vector(31 downto 0);5��    
                     �                      �    
                     �                      �    
                     �                      �                         �                      �                         �                      5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                                                V       e��H     �         D      :    signal q_expected, q_actual : bit_vector(31 downto 0);5��              	           �       	               5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                                                V       e��K     �         D      1    signal q, q_actual : bit_vector(31 downto 0);5��                         �                      5�_�   4   8           5          ����                                                                                                                                                                                                                                                                                                                                                V       e��S     �         D      &    signal q: bit_vector(31 downto 0);5��                         �                      5�_�   5   9   6       8          ����                                                                                                                                                                                                                                                                                                                                                V       e��b     �         D      E        port map (x => x_tb, y => y_tb, z => z_tb, q => q_tb_actual);5��                        %                    5�_�   8   :           9          ����                                                                                                                                                                                                                                                                                                                                                V       e��e    �         D      B        port map (x => x, y => y_tb, z => z_tb, q => q_tb_actual);5��                        -                    5�_�   9   ;           :      '    ����                                                                                                                                                                                                                                                                                                                                                V       e��h     �         D      ?        port map (x => x, y => y, z => z_tb, q => q_tb_actual);5��       '                 5                    5�_�   :   <           ;      /    ����                                                                                                                                                                                                                                                                                                                                                V       e��l     �         D      <        port map (x => x, y => y, z => z, q => q_tb_actual);5��       /                 =                    5�_�   ;   =           <   
        ����                                                                                                                                                                                                                                                                                                                            
   	                  V   	    e��{     �   
                  -- Signals for the testbench   -    signal x, y, z : bit_vector(31 downto 0);   '    signal q : bit_vector(31 downto 0);    �   	   
   H           -- Signals for the testbench   -    signal x, y, z : bit_vector(31 downto 0);   '    signal q : bit_vector(31 downto 0);    �         D    5��   	              
       �       x       �       5�_�   <   >           =           ����                                                                                                                                                                                                                                                                                                                               	                  V   	    e��|     �                     -- Signals for the testbench   -    signal x, y, z : bit_vector(31 downto 0);   '    signal q : bit_vector(31 downto 0);    �   
      H           -- Signals for the testbench   -    signal x, y, z : bit_vector(31 downto 0);   '    signal q : bit_vector(31 downto 0);    �         D    5��   
                     �       x       �       �                                              �                         2                    5�_�   =   ?           >           ����                                                                                                                                                                                                                                                                                                                               	                  V   	    e��|     �                     -- Signals for the testbench   1        signal x, y, z : bit_vector(31 downto 0);   +        signal q : bit_vector(31 downto 0);    �         H           -- Signals for the testbench   1        signal x, y, z : bit_vector(31 downto 0);   +        signal q : bit_vector(31 downto 0);    �         D    5��                        �       �       �       �                         �                     5�_�   >   @           ?           ����                                                                                                                                                                                                                                                                                                                               	                  V   	    e��|     �                $        -- Signals for the testbench   1        signal x, y, z : bit_vector(31 downto 0);   +        signal q : bit_vector(31 downto 0);    �         H      $        -- Signals for the testbench   1        signal x, y, z : bit_vector(31 downto 0);   +        signal q : bit_vector(31 downto 0);    �         D    5��                        �       �             5�_�   ?   A           @           ����                                                                                                                                                                                                                                                                                                                               	                  V   	    e��|     �                $        -- Signals for the testbench   1        signal x, y, z : bit_vector(31 downto 0);   +        signal q : bit_vector(31 downto 0);    �         H      $        -- Signals for the testbench   1        signal x, y, z : bit_vector(31 downto 0);   +        signal q : bit_vector(31 downto 0);    �         D    5��                              �       J      �                         o                    5�_�   @   B           A           ����                                                                                                                                                                                                                                                                                                                               	                  V   	    e��}     �                $        -- Signals for the testbench   5            signal x, y, z : bit_vector(31 downto 0);   +        signal q : bit_vector(31 downto 0);    �         H      $        -- Signals for the testbench   5            signal x, y, z : bit_vector(31 downto 0);   +        signal q : bit_vector(31 downto 0);    �         D    5��                        J      �       U      �                         U                    �                         ~                    5�_�   A   C           B           ����                                                                                                                                                                                                                                                                                                                               	                  V   	    e��}     �                (            -- Signals for the testbench   1        signal x, y, z : bit_vector(31 downto 0);   +        signal q : bit_vector(31 downto 0);    �         H      (            -- Signals for the testbench   1        signal x, y, z : bit_vector(31 downto 0);   +        signal q : bit_vector(31 downto 0);    �         D    5��                        U      �       h      �                         h                    �                         �                    �                         �                    5�_�   B   D           C           ����                                                                                                                                                                                                                                                                                                                               	                  V   	    e��}     �                $        -- Signals for the testbench   -    signal x, y, z : bit_vector(31 downto 0);   '    signal q : bit_vector(31 downto 0);    �         H      $        -- Signals for the testbench   -    signal x, y, z : bit_vector(31 downto 0);   '    signal q : bit_vector(31 downto 0);    �         D    5��                        h      |       i      �                         i                    5�_�   C   E           D          ����                                                                                                                                                                                                                                                                                                                               	                  V   	    e�ނ     �         D      '    signal q : bit_vector(31 downto 0);5��                        �                    5�_�   D   H           E      /    ����                                                                                                                                                                                                                                                                                                                               	                  V   	    e�އ     �         D      2        port map (x => x, y => y, z => z, q => q);5��       /                 A                    5�_�   E   I   F       H           ����                                                                                                                                                                                                                                                                                                                                      	           V       e���    �                    -- Constants   (    constant CLK_PERIOD : time := 10 ns;    5��                          V       ;               5�_�   H   J           I   *       ����                                                                                                                                                                                                                                                                                                                                                 V       e��%     �   *   ,   B              �   *   ,   A    5��    *                      I              	       �    *                     Q                     �    *                     I                    �    *                     Q                     �    *   
                 S                    5�_�   I   K           J   +       ����                                                                                                                                                                                                                                                                                                                                                 V       e��+     �   *   +              end loop;5��    *                      I                     5�_�   J   L           K   (        ����                                                                                                                                                                                                                                                                                                                                       (           V       e��6     �      )   A   	   '        while not endfile(tb_file) loop               -- read inputs   '            readline(tb_file, tb_line);               read(tb_line, Xv);               X <= signed(Xv);   !            read(tb_line, space);               read(tb_line, Bv);               B <= signed(Bv);    5��           	       	                    (      5�_�   K   M           L   ,        ����                                                                                                                                                                                                                                                                                                                            ,           =           V        e��D     �   +   ,                  -- Check results process   "    check_results_process: process   	    begin   '        for i in test_vector'range loop   7            -- Allow time for the DUT to produce output                wait for CLK_PERIOD;       B            -- Apply the expected output for the current test case   -            q_tb_expected <= (others => '0');   .            assert q_tb_actual = q_tb_expected   F                report "Test case " & integer'image(i + 1) & " failed"   !                severity failure;       K            -- Add more result checking as needed for the current test case           end loop;               wait;5��    +                      |      D              5�_�   L   N           M   ,        ����                                                                                                                                                                                                                                                                                                                            ,           ,           V        e��E     �   +   ,              end process;5��    +                      |                     5�_�   M   O           N   ,        ����                                                                                                                                                                                                                                                                                                                            ,           ,           V        e��F     �   +   ,           5��    +                      |                     5�_�   N   P           O   (        ����                                                                                                                                                                                                                                                                                                                            ,           ,           V        e��V     �   '   )   -      
        --5��    '                    %                    �    '                     (                     �    '   
                  '                     �    '   	                  &                     �    '                    %                    �    '                    %                    �    '                    %                    �    '                 2   %             2       5�_�   O   Q           P   (       ����                                                                                                                                                                                                                                                                                                                            (          (          v       e��Y     �   '   )   -      :        assert neg_condition report message severity note;5��    '                    ,                    5�_�   P   R           Q   (       ����                                                                                                                                                                                                                                                                                                                            (   "       (          v       e��[     �   '   )   -      2        assert false report message severity note;5��    '                     9                     5�_�   Q   S           R   (       ����                                                                                                                                                                                                                                                                                                                            (   "       (          v       e��[     �   '   )   -      +        assert false report  severity note;5��    '                     9                     5�_�   R   T           S   (       ����                                                                                                                                                                                                                                                                                                                            (   "       (          v       e��[    �   '   )   -      -        assert false report "" severity note;5��    '                     :                     5�_�   S   U           T   (   )    ����                                                                                                                                                                                                                                                                                                                            (   )       (   )       V   )    e�߰     �   '   (          0        assert false report "BOT" severity note;5��    '                            1               5�_�   T   V           U            ����                                                                                                                                                                                                                                                                                                                            (   )       (   )       V   )    e�߲     �      !   ,    �       !   ,    5��                                         1       5�_�   U   W           V           ����                                                                                                                                                                                                                                                                                                                            )   )       )   )       V   )    e�߲     �       "   -    5��                           1              	       �                          8                     �                          7                     �                          6                     �                          5                     �                          4                     �                          3                     �                          2                     �                           1                     5�_�   V   X           W            ����                                                                                                                                                                                                                                                                                                                            *   )       *   )       V   )    e�ߴ    �      !   /              �      !   .    5��                                         	       �                                              5�_�   W   Y           X   !        ����                                                                                                                                                                                                                                                                                                                            +   )       +   )       V   )    e��    �       "   /      0        assert false report "BOT" severity note;5��                           <                     �        !                 =                    5�_�   X   Z           Y   !        ����                                                                                                                                                                                                                                                                                                                            +   )       +   )       V   )    e��.     �       "   /      8        assert false report "BOT \n baba" severity note;5��                           <                     5�_�   Y   [           Z   !   !    ����                                                                                                                                                                                                                                                                                                                            +   )       +   )       V   )    e��1     �       "   /      0        assert false report "BOT" severity note;5��        !                  =                     �        %                 A                    5�_�   Z   \           [   !   +    ����                                                                                                                                                                                                                                                                                                                            +   )       +   )       V   )    e��;     �       "   /      :        assert false report "BOT" & x'image severity note;5��        +                  G                     5�_�   [   ]           \   !   ,    ����                                                                                                                                                                                                                                                                                                                            +   )       +   )       V   )    e��@     �       "   /      <        assert false report "BOT" & x'image() severity note;5��        ,                  H                     5�_�   \   ^           ]   !   $    ����                                                                                                                                                                                                                                                                                                                            +   )       +   )       V   )    e��B     �       "   /      =        assert false report "BOT" & x'image(x) severity note;5��        $                 @                    5�_�   ]   `           ^   !   $    ����                                                                                                                                                                                                                                                                                                                            +   )       +   )       V   )    e��L     �       "   /      C        assert false report "BOT" & integer'image(x) severity note;5��        $                 @                    �        &                  B                     �        %                  A                     �        $              
   @             
       �        $       
          @      
              �        $              
   @             
       5�_�   ^   a   _       `           ����                                                                                                                                                                                                                                                                                                                            +   )       +   )       V   )    e���     �         /    �         /    5��                          �              ,       5�_�   `   b           a          ����                                                                                                                                                                                                                                                                                                                            ,   )       ,   )       V   )    e���     �         0      +    signal saida : bit_vector(31 downto 0);5��                         �                     5�_�   a   d           b          ����                                                                                                                                                                                                                                                                                                                            ,   )       ,   )       V   )    e���    �         0      ,    signal saidai : bit_vector(31 downto 0);5��                        �                    5�_�   b   e   c       d          ����                                                                                                                                                                                                                                                                                                                            ,   )       ,   )       V   )    e���     �         1          �         1    �         0    5��                          �                     �                       *   �              *       �       *                 �                     �                          �                     5�_�   d   f           e          ����                                                                                                                                                                                                                                                                                                                            .   )       .   )       V   )    e��    �         2          signal saidai : integer;5��                         �                     �                        �                    �       '                 �                    5�_�   e   g           f   $   $    ����                                                                                                                                                                                                                                                                                                                            .   )       .   )       V   )    e��$     �   #   %   2      F        assert false report "BOT" & bit_vector'image(x) severity note;5��    #   $       
          �      
              5�_�   f   h           g   $   2    ����                                                                                                                                                                                                                                                                                                                            .   )       .   )       V   )    e��(    �   #   %   2      C        assert false report "BOT" & integer'image(x) severity note;5��    #   2                 �                    �    #   4                  �                     �    #   3                  �                     �    #   2                 �                    �    #   6                  �                     �    #   5                  �                     �    #   4                  �                     �    #   3                  �                     �    #   2                 �                    �    #   3                  �                     �    #   2                 �                    �    #   2                 �                    �    #   2                 �                    5�_�   g   j           h          ����                                                                                                                                                                                                                                                                                                                            .   )       .   )       V   )    e��X    �         3       �         3    �         2    5��                          "                      �                         "               P       5�_�   h   k   i       j          ����                                                                                                                                                                                                                                                                                                                            1   )       1   )       V   )    e��h     �                use ieee.numeric_std.ALL;5��                          Y                      5�_�   j   l           k           ����                                                                                                                                                                                                                                                                                                                            0   )       0   )       V   )    e��j    �                use ieee.std_logic_1164.ALL;5��                          "                      5�_�   k   m           l   /        ����                                                                                                                                                                                                                                                                                                                            /   )       /   )       V   )    e���     �   /   1   3    �   /   0   3    5��    /                      �              I       5�_�   l   n           m   0       ����                                                                                                                                                                                                                                                                                                                            /   )       /   )       V   )    e���     �   /   1   4      H        assert false report "BOT" & integer'image(saidai) severity note;5��    /                                        5�_�   m   o           n   0   "    ����                                                                                                                                                                                                                                                                                                                            /   )       /   )       V   )    e���     �   /   1   4      H        assert false report "EOT" & integer'image(saidai) severity note;5��    /   "                                       5�_�   n   p           o   0   "    ����                                                                                                                                                                                                                                                                                                                            /   )       /   )       V   )    e���    �   /   1   4      8        assert false report "EOT" saidai) severity note;5��    /   "                                       5�_�   o   q           p   %        ����                                                                                                                                                                                                                                                                                                                            /   )       /   )       V   )    e��'     �   $   &   4      H        assert false report "BOT" & integer'image(saidai) severity note;5��    $                      �                     5�_�   p   r           q   %   #    ����                                                                                                                                                                                                                                                                                                                            /   )       /   )       V   )    e��.     �   $   &   4      K        assert false report "BOT ch" & integer'image(saidai) severity note;5��    $   #               	   �              	       5�_�   q   t           r   0        ����                                                                                                                                                                                                                                                                                                                            /   )       /   )       V   )    e��3    �   /   1   4      0        assert false report "EOT" severity note;5��    /                      !                     5�_�   r   u   s       t   .       ����                                                                                                                                                                                                                                                                                                                            '          .          V       e��}     �   &   /   4      *        -- while not endfile(tb_file) loop           --     -- read inputs   *        --     readline(tb_file, tb_line);   !        --     read(tb_line, Xv);           --     X <= signed(Xv);   $        --     read(tb_line, space);   !        --     read(tb_line, Bv);           --     B <= signed(Bv);5��    &                     �                  5�_�   t   v           u   '        ����                                                                                                                                                                                                                                                                                                                            '          /           V       e��     �   &   '       	   '        while not endfile(tb_file) loop               -- read inputs   '            readline(tb_file, tb_line);               read(tb_line, Xv);               X <= signed(Xv);   !            read(tb_line, space);               read(tb_line, Bv);               B <= signed(Bv);    5��    &       	               �                    5�_�   u   w           v   "        ����                                                                                                                                                                                                                                                                                                                            '          '           V       e��     �   "   ,   +    �   "   #   +    5��    "               	       g                    5�_�   v   x           w   *       ����                                                                                                                                                                                                                                                                                                                            0          0           V       e��O     �   *   ,   5                  �   *   ,   4    5��    *                      l                     �    *                     x                     �    *                     l                    �    *                     x                     5�_�   w   y           x   "        ����                                                                                                                                                                                                                                                                                                                            +          "           V       e��p     �   !   "       
       '        while not endfile(tb_file) loop               -- read inputs   '            readline(tb_file, tb_line);               read(tb_line, Xv);               X <= signed(Xv);   !            read(tb_line, space);               read(tb_line, Bv);               B <= signed(Bv);           end loop;5��    !       
               f                    5�_�   x   z           y   $        ����                                                                                                                                                                                                                                                                                                                            "          "           V       e��r     �   $   /   +    �   $   %   +    5��    $               
       �                    5�_�   y   {           z   .        ����                                                                                                                                                                                                                                                                                                                            "          "           V       e��u     �   .   0   5    5��    .                      �              	       �    .                      �                     5�_�   z   |           {   *       ����                                                                                                                                                                                                                                                                                                                            "          "           V       e���     �   )   +   6                  X <= signed(Xv);5��    )                     )                     5�_�   {   }           |   *       ����                                                                                                                                                                                                                                                                                                                            "          "           V       e���     �   )   +   6                  X <= (Xv);5��    )                     )                     5�_�   |   ~           }   *       ����                                                                                                                                                                                                                                                                                                                            "          "           V       e���     �   )   +   6                  X <= Xv);5��    )                     +                     5�_�   }              ~   !       ����                                                                                                                                                                                                                                                                                                                            "          "           V       e���     �       "   6      :        variable Xv, Yv, Zv, res: bit_vector(31 downto 0);5��                          +      ;       >       5�_�   ~   �              )       ����                                                                                                                                                                                                                                                                                                                            "          "           V       e���     �   (   *   6                  read(tb_line, Xv);5��    (                                        5�_�      �           �   *       ����                                                                                                                                                                                                                                                                                                                            "          "           V       e���     �   )   *                      X <= Xv;5��    )                                           5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            "          "           V       e���     �   *   ,   5                  read(tb_line, Bv);5��    *                    V                    5�_�   �   �           �   +        ����                                                                                                                                                                                                                                                                                                                            *          +          V       e��      �   +   .   5    �   +   ,   5    5��    +                      Z              @       5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                            *          +          V       e��     �   ,   .   7                  read(tb_line, y);5��    ,                    �                    5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            *          +          V       e��     �   -   .                      B <= signed(Bv);5��    -                      �                     5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                            *          +          V       e��     �   (   *   6    5��    (                      �                     �    (                      �                     5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            +          ,          V       e��     �   .   0   7    5��    .                      �                     �    .                      �                     5�_�   �   �           �   .        ����                                                                                                                                                                                                                                                                                                                            +          ,          V       e��c     �   .   0   8    �   .   /   8    5��    .                      �              U       5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            +          ,          V       e��d     �   .   0   9      T        assert false report "BOT ch function" & integer'image(saidai) severity note;5��    .                     �                     5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            +          ,          V       e��f     �   .   0   9    5��    .                      �                     �    .                      �                     5�_�   �   �           �   0   !    ����                                                                                                                                                                                                                                                                                                                            +          ,          V       e��k     �   /   1   :      X            assert false report "BOT ch function" & integer'image(saidai) severity note;5��    /   !                 �                    5�_�   �   �           �   0   8    ����                                                                                                                                                                                                                                                                                                                            +          ,          V       e��     �   /   1   :      N            assert false report "x is " & integer'image(saidai) severity note;5��    /   8                 �                    �    /   9                  �                     �    /   8              
   �             
       �    /   8       
          �      
              �    /   8              
   �             
       5�_�   �   �           �   0   B    ����                                                                                                                                                                                                                                                                                                                            +          ,          V       e��     �   /   1   :      R            assert false report "x is " & integer'image(to_integer) severity note;5��    /   B                  �                     5�_�   �   �           �   0   C    ����                                                                                                                                                                                                                                                                                                                            +          ,          V       e��     �   /   1   :      T            assert false report "x is " & integer'image(to_integer()) severity note;5��    /   C                  �                     �    /   E                  �                     �    /   D                  �                     �    /   C                 �                    �    /   J                  �                     �    /   I                  �                     �    /   H                  �                     �    /   G                  �                     �    /   F                  �                     �    /   E                  �                     �    /   D                  �                     �    /   C                 �                    �    /   E                  �                     �    /   D                  �                     �    /   C                 �                    �    /   J                  �                     �    /   I                  �                     �    /   H                  �                     �    /   G                  �                     �    /   F                  �                     �    /   E                  �                     �    /   D                  �                     �    /   C                 �                    �    /   E                  �                     �    /   D                  �                     �    /   C                 �                    �    /   J                  �                     �    /   I                  �                     �    /   H                  �                     �    /   G                  �                     �    /   F                  �                     �    /   E                  �                     �    /   D                  �                     �    /   C                 �                    �    /   C                 �                    �    /   C              	   �             	       �    /   K                  �                     5�_�   �   �           �   0   K    ����                                                                                                                                                                                                                                                                                                                            +          ,          V       e��     �   /   1   :      \            assert false report "x is " & integer'image(to_integer(unsigned)) severity note;5��    /   K                  �                     5�_�   �   �           �   0   L    ����                                                                                                                                                                                                                                                                                                                            +          ,          V       e��     �   /   1   :      ^            assert false report "x is " & integer'image(to_integer(unsigned())) severity note;5��    /   L                  �                     5�_�   �   �           �   0   C    ����                                                                                                                                                                                                                                                                                                                            +          ,          V       e��    �   /   1   :      _            assert false report "x is " & integer'image(to_integer(unsigned(x))) severity note;5��    /   C                 �                    5�_�   �   �           �   !   <    ����                                                                                                                                                                                                                                                                                                                            +          ,          V       e��     �       "   :      =        -- variable Xv, Yv, Zv, res: bit_vector(31 downto 0);5��                          +      >       ;       5�_�   �   �           �   *       ����                                                                                                                                                                                                                                                                                                                            +          ,          V       e��     �   *   ,   ;                  �   *   ,   :    5��    *                                           �    *                     $                     5�_�   �   �           �   *       ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e���     �   )   +   ;                  read(tb_line, x);5��    )                                        5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��     �   -   /   ;    �   -   .   ;    5��    -                      n                     5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��     �   ,   .   <                  read(tb_line, y);5��    ,                    j                    5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��	     �   -   /   <                  x <= Xv;5��    -                    �                    5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��
     �   -   /   <                  x <= Yv;5��    -                    {                    5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��     �   /   1   <                  read(tb_line, z);5��    /                    �                    5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��     �   0   2   <    �   0   1   <    5��    0                      �                     5�_�   �   �           �   1       ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��     �   0   2   =                  y <= Yv;5��    0                    �                    5�_�   �   �           �   1       ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��    �   0   2   =                  z <= Yv;5��    0                    �                    5�_�   �   �           �   3   C    ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��V    �   2   4   =      ]            assert false report "x is " & integer'image(to_integer(signed(x))) severity note;5��    2   C                                     �    2   E                                        �    2   D                                       �    2   C                                     �    2   E                                        �    2   D                                       �    2   C                                     �    2   C                                     �    2   C                                     �    2   C                                     5�_�   �   �           �   3   M    ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��   " �   2   4   =      _            assert false report "x is " & integer'image(to_integer(unsigned(x))) severity note;5��    2   L                 '                    5�_�   �   �   �       �   3   C    ����                                                                                                                                                                                                                                                                                                                                                             e�
]   # �   2   4   =      `            assert false report "x is " & integer'image(to_integer(unsigned(Xv))) severity note;5��    2   C                                     5�_�   �   �           �   1       ����                                                                                                                                                                                                                                                                                                                                                             e�
|     �   1   4   >                  �   1   3   =    5��    1                      �                     �    1                      �                     �    1                     �                     �    2                  	   �              	       5�_�   �   �           �   3       ����                                                                                                                                                                                                                                                                                                                                                             e�
�     �   2   4   ?                  wait 1ns;5��    2                     �                     5�_�   �   �           �   3       ����                                                                                                                                                                                                                                                                                                                                                             e�
�     �   2   4   ?                  wait 1 ns;5��    2                     �                     5�_�   �   �           �   5   J    ����                                                                                                                                                                                                                                                                                                                                                             e�
�   $ �   4   6   ?      ^            assert false report "x is " & integer'image(to_integer(signed(Xv))) severity note;5��    4   J                 A                    5�_�   �   �           �   5   J    ����                                                                                                                                                                                                                                                                                                                                                             e�
�     �   5   7   @                  �   5   7   ?    5��    5                      U                     �    5                     a                     �    5                     c                     �    5                     b                     �    5                    a                    �    5                    a                    �    5                    a                    �    5                 2   a             2       5�_�   �   �           �   6       ����                                                                                                                                                                                                                                                                                                                            6          6          v       e�     �   5   7   @      >            assert neg_condition report message severity note;5��    5                    h                    �    5                     m                     5�_�   �   �           �   6        ����                                                                                                                                                                                                                                                                                                                            6   &       6           v        e�     �   5   7   @      6            assert x = y report message severity note;5��    5                      u                     5�_�   �   �           �   6        ����                                                                                                                                                                                                                                                                                                                            6   &       6           v        e�     �   5   7   @      /            assert x = y report  severity note;5��    5                      u                     5�_�   �   �           �   6   !    ����                                                                                                                                                                                                                                                                                                                            6   &       6           v        e�     �   5   7   @      1            assert x = y report "" severity note;5��    5   !               
   v              
       5�_�   �   �           �   6       ����                                                                                                                                                                                                                                                                                                                            6   &       6           v        e�   % �   5   7   @      ;            assert x = y report "x equals y" severity note;5��    5                     j                     �    5                    j                    5�_�   �   �           �   :       ����                                                                                                                                                                                                                                                                                                                            6   &       6           v        e�h     �   9   :          T        assert false report "BOT ch function" & integer'image(saidai) severity note;5��    9                      �      U               5�_�   �   �           �   $        ����                                                                                                                                                                                                                                                                                                                            6   &       6           v        e�j     �   $   &   ?    �   $   %   ?    5��    $                      �              U       5�_�   �   �           �   <       ����                                                                                                                                                                                                                                                                                                                            7   &       7           v        e�m     �   <   >   @    5��    <                      9              	       �    <                     @                     �    <                     ?                     �    <                     >                     �    <                     =                     �    <                     <                     �    <                     ;                     �    <                     :                     �    <                      9                     5�_�   �   �           �   <        ����                                                                                                                                                                                                                                                                                                                            7   &       7           v        e�o     �   ;   =   B              �   ;   =   A    5��    ;                      �              	       �    ;                                          5�_�   �   �           �   ;        ����                                                                                                                                                                                                                                                                                                                            7   &       7           v        e�t     �   :   ;           5��    :                      �                     5�_�   �   �           �   4       ����                                                                                                                                                                                                                                                                                                                            7   &       7           v        e�|     �   4   7   B                  �   4   6   A    5��    4                      K                     �    4                      K                     �    4                     K                     �    5                     W                     �    5   
                  V                     �    5   	                  U                     �    5                     T                     �    5                     S                     �    5                     R                     �    5                     Q                     �    5                     P                     �    5                     O                     �    5                     N                     �    5                     M                     �    5                      L                     5�_�   �   �           �   6        ����                                                                                                                                                                                                                                                                                                                            9   &       9           v        e��     �   5   6               5��    5                      L                     5�_�   �   �           �   6   !    ����                                                                                                                                                                                                                                                                                                                            7   &       7           v        e��     �   5   7   A      ]            assert false report "x is " & integer'image(to_integer(signed(x))) severity note;5��    5   !                 m                    5�_�   �   �           �   6   "    ����                                                                                                                                                                                                                                                                                                                            7   &       7           v        e��     �   5   7   A      ]            assert false report "F is " & integer'image(to_integer(signed(x))) severity note;5��    5   !                 m                    5�_�   �   �           �   6   O    ����                                                                                                                                                                                                                                                                                                                            7   &       7           v        e��   & �   5   7   A      b            assert false report "output is " & integer'image(to_integer(signed(x))) severity note;5��    5   O                 �                    5�_�   �   �           �   6   P    ����                                                                                                                                                                                                                                                                                                                            7   &       7           v        e��   ' �   5   7   A      b            assert false report "output is " & integer'image(to_integer(signed(q))) severity note;5��    5   O                 �                    5�_�   �   �           �   2        ����                                                                                                                                                                                                                                                                                                                            0           2          V   S    e��     �   2   6   A    �   2   3   A    5��    2                      /              V       5�_�   �   �           �   4       ����                                                                                                                                                                                                                                                                                                                            0           2          V   S    e�    ( �   3   5   D                  read(tb_line, Zv);5��    3                    k                    5�_�   �   �           �   5       ����                                                                                                                                                                                                                                                                                                                            0           2          V   S    e�%   ) �   4   5                      z <= Zv;5��    4                      q                     5�_�   �   �           �   8        ����                                                                                                                                                                                                                                                                                                                            0           2          V   S    e�0     �   8   :   C    �   8   9   C    5��    8                      �              g       5�_�   �   �           �   9   !    ����                                                                                                                                                                                                                                                                                                                            0           2          V   S    e�3     �   8   :   D      f            assert false report "output is " & integer'image(to_integer(signed(saida))) severity note;5��    8   !               	                 	       5�_�   �   �           �   9   X    ����                                                                                                                                                                                                                                                                                                                            0           2          V   S    e�:   * �   8   :   D      o            assert false report "expected output is " & integer'image(to_integer(signed(saida))) severity note;5��    8   X                 M                    5�_�   �   �           �   %   .    ����                                                                                                                                                                                                                                                                                                                            %   D       %   .       v   .    e�o     �   $   &   D      T        assert false report "BOT ch function" & integer'image(saidai) severity note;5��    $   .                  �                     5�_�   �   �           �   %   -    ����                                                                                                                                                                                                                                                                                                                            %   D       %   .       v   .    e�q   + �   $   &   D      =        assert false report "BOT ch function"  severity note;5��    $   -                  �                     5�_�   �   �           �   9   -    ����                                                                                                                                                                                                                                                                                                                            %   D       %   .       v   .    e�)�     �   9   ;   E                  �   9   ;   D    5��    9                      K                     �    9                     W                     �    9                     Y                     �    9                     X                     �    9                    W                    �    9                    W                    �    9                    W                    �    9                 2   W             2       5�_�   �   �           �   :       ����                                                                                                                                                                                                                                                                                                                            :          :          v       e�)�     �   9   ;   E      >            assert neg_condition report message severity note;5��    9                    ^                    �    9                     _                     �    9                    ^                    �    9                    ^                    �    9                    ^                    �    9                     i                     5�_�   �   �           �   :   &    ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�)�     �   9   ;   E      <            assert saida = res report message severity note;5��    9   &                  q                     5�_�   �   �           �   :   &    ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�)�     �   9   ;   E      5            assert saida = res report  severity note;5��    9   &                  q                     5�_�   �   �           �   :   '    ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�)�     �   9   <   E      7            assert saida = res report "" severity note;5��    9   '                  r                     �    9   (                  s                     �    9   '                  r                     �    9   &                  q                     �    9   &                  q                     �    9   %                  p                     �    9   %                p                    5�_�   �   �           �   ;       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�)�     �   :   <   F    5��    :                      q                     5�_�   �   �           �   ;       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�)�     �   :   <   G                  5��    :                     }                     5�_�   �   �           �   ;       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�)�     �   :   <   G                  ""5��    :                     ~                     5�_�   �   �           �   ;       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�)�     �   :   =   G                  "Output failed"5��    :                     �                     �    :                    �                     5�_�   �   �           �   <       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*     �   ;   =   H                  5��    ;                     �                     5�_�   �   �           �   <       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*)   , �   ;   =   H                  ""5��    ;                     �                     5�_�   �   �           �   =       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*1   - �   <   >   H                  severity note;5��    <                    �                    5�_�   �   �           �   ;       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*A   . �   :   <   H                  "Output failed" &5��    :                     �                     �    :                    �                    5�_�   �   �           �   <       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*Z     �   ;   =   H                  "trst"5��    ;                     �                     �    ;                     �                     �    ;                     �                     �    ;                    �                    �    ;                    �                    �    ;                     �                     �    ;                     �                     �    ;                    �                    5�_�   �   �           �   <       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*f     �   ;   =   H                  " X="5��    ;                     �                     �    ;                     �                     �    ;                    �                    �    ;                     �                     �    ;                     �                     �    ;                     �                     �    ;                    �                    �    ;                     �                     �    ;                     �                     �    ;                     �                     �    ;                     �                     �    ;                     �                     �    ;                     �                     �    ;                    �                    �    ;                    �                    �    ;                 
   �             
       �    ;                     �                     �    ;                    �                    �    ;                    �                    �    ;                    �                    5�_�   �   �           �   <   !    ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*x     �   ;   =   H      !            " X=" & integer'image5��    ;   !                  �                     5�_�   �   �           �   <   "    ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*y     �   ;   =   H      #            " X=" & integer'image()5��    ;   "                  �                     �    ;   #                  �                     �    ;   "              
   �             
       �    ;   "       
          �      
              �    ;   "              
   �             
       5�_�   �   �           �   <   ,    ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*{     �   ;   =   H      -            " X=" & integer'image(to_integer)5��    ;   ,                  �                     5�_�   �   �           �   <   -    ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*|     �   ;   =   H      /            " X=" & integer'image(to_integer())5��    ;   -                  �                     �    ;   /                  �                     �    ;   .                  �                     �    ;   -                 �                    �    ;   -                 �                    �    ;   -                 �                    5�_�   �   �           �   <   3    ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*~     �   ;   =   H      5            " X=" & integer'image(to_integer(signed))5��    ;   3                  �                     5�_�   �   �           �   <   4    ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*     �   ;   =   H      7            " X=" & integer'image(to_integer(signed()))5��    ;   4                  �                     5�_�   �   �           �   <   4    ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*�     �   <   >   H    �   <   =   H    5��    <                      �              9       5�_�   �   �           �   =       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*�     �   =   ?   I    �   =   >   I    5��    =                                    9       5�_�   �   �           �   =       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*�     �   <   >   J      8            " X=" & integer'image(to_integer(signed(x)))5��    <                    �                    5�_�   �   �           �   =   4    ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*�     �   <   >   J      8            " Y=" & integer'image(to_integer(signed(x)))5��    <   4                 �                    5�_�   �   �           �   >   4    ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*�     �   =   ?   J      8            " X=" & integer'image(to_integer(signed(x)))5��    =   4                 8                    5�_�   �   �           �   >       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*�     �   =   ?   J      8            " X=" & integer'image(to_integer(signed(z)))5��    =                                        5�_�   �   �           �   >       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*�     �   =   ?   J      8            " |=" & integer'image(to_integer(signed(z)))5��    =                                        5�_�   �   �           �   >       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*�     �   >   @   J    �   >   ?   J    5��    >                      =              9       5�_�   �   �           �   ?       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*�     �   ?   A   K    �   ?   @   K    5��    ?                      v              9       5�_�   �   �           �   ?       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*�     �   >   @   L      8            " X=" & integer'image(to_integer(signed(x)))5��    >                 
   K             
       5�_�   �   �           �   @       ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*�     �   ?   A   L      8            " X=" & integer'image(to_integer(signed(x)))5��    ?                 
   �             
       5�_�   �   �           �   ?   >    ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*�     �   >   @   L      A            " Computed Q=" & integer'image(to_integer(signed(x)))5��    >   =                 z                    5�_�   �   �           �   @   =    ����                                                                                                                                                                                                                                                                                                                            :   ,       :   &       v   &    e�*�     �   ?   A   L      A            " Expected Q=" & integer'image(to_integer(signed(x)))5��    ?   =                 �                    5�_�   �   �           �   <   8    ����                                                                                                                                                                                                                                                                                                                            <   7       >   8          ?    e�*�     �   <   ?   L      8            " Y=" & integer'image(to_integer(signed(y)))   8            " Z=" & integer'image(to_integer(signed(z)))�   ;   =   L      8            " X=" & integer'image(to_integer(signed(x)))5��    ;   8                  �                     �    <   8                                       �    =   8                  F                     5�_�   �   �           �   ?   E    ����                                                                                                                                                                                                                                                                                                                            <   7       >   8          ?    e�*�     �   >   @   L      E            " Computed Q=" & integer'image(to_integer(signed(saida)))5��    >   E                  �                     5�_�   �   �           �   B   ;    ����                                                                                                                                                                                                                                                                                                                            <   7       >   8          ?    e�*�     �   A   B          <            assert x /= y report "x equals y" severity note;5��    A                      �      =               5�_�   �   �           �   8        ����                                                                                                                                                                                                                                                                                                                            <   7       >   8          ?    e�*�   / �   7   8          f            assert false report "output is " & integer'image(to_integer(signed(saida))) severity note;   m            assert false report "expected output is " & integer'image(to_integer(signed(res))) severity note;5��    7                      v      �               5�_�   �   �           �   8       ����                                                                                                                                                                                                                                                                                                                            :   7       <   8          ?    e�7�     �   7   9   I      %            assert saida = res report5��    7                    �                    5�_�   �   �           �   8       ����                                                                                                                                                                                                                                                                                                                            :   7       <   8          ?    e�7�     �   7   9   I      &            assert signed = res report5��    7                     �                     5�_�   �   �           �   8       ����                                                                                                                                                                                                                                                                                                                            :   7       <   8          ?    e�7�     �   7   9   I      (            assert signed() = res report�   8   9   I    5��    7                     �                     5�_�   �   �           �   8   #    ����                                                                                                                                                                                                                                                                                                                            :   7       <   8          ?    e�7�     �   7   9   I      -            assert signed(saida) = res report5��    7   #                 �                    5�_�   �   �           �   8   )    ����                                                                                                                                                                                                                                                                                                                            :   7       <   8          ?    e�7�     �   7   9   I      0            assert signed(saida) = signed report5��    7   )                  �                     5�_�   �   �           �   8   )    ����                                                                                                                                                                                                                                                                                                                            :   7       <   8          ?    e�7�   0 �   7   9   I      2            assert signed(saida) = signed() report�   8   9   I    5��    7   *                  �                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            :   7       <   8          ?    e�7�   1 �         I      *    saidai <= to_integer(unsigned(saida));5��                                            5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            :   7       <   8          ?    e�7�     �                (    saidai <= to_integer(signed(saida));5��                          �      )               5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            9   7       ;   8          ?    e�7�   2 �                *    signal saidai : integer range 0 to 31;5��                          �      +               5�_�   �   �           �   6       ����                                                                                                                                                                                                                                                                                                                            8   7       :   8          ?    e�7�     �   5   7   G      5            assert signed(saida) = signed(res) report5��    5                     3                     5�_�   �   �           �   6       ����                                                                                                                                                                                                                                                                                                                            8   7       :   8          ?    e�7�     �   5   7   G      /            assert (saida) = signed(res) report5��    5                     3                     5�_�   �   �           �   6       ����                                                                                                                                                                                                                                                                                                                            8   7       :   8          ?    e�7�     �   5   7   G      .            assert saida) = signed(res) report5��    5                     8                     5�_�   �              �   6       ����                                                                                                                                                                                                                                                                                                                            8   7       :   8          ?    e�7�     �   5   7   G      -            assert saida = signed(res) report5��    5                     ;                     5�_�   �                6       ����                                                                                                                                                                                                                                                                                                                            8   7       :   8          ?    e�7�   3 �   5   7   G      &            assert saida = res) report5��    5                     >                     5�_�                     4    ����                                                                                                                                                                                                                                                                                                                            8   7       :   8          ?    e�9i   4 �         G      :        file tb_file : text open read_mode is "cases.dat";5��       4                  �                     5�_�                  /    ����                                                                                                                                                                                                                                                                                                                                       G           V        e�<�     �         G      =        file tb_file : text open read_mode is "cases_ch.dat";5��       /                  �                     �       /                  �                     5�_�                    /    ����                                                                                                                                                                                                                                                                                                                                       G           V        e�<�   9 �         G      =        file tb_file : text open read_mode is "cases_ch.dat";5��       /                 �                    5�_�               8       ����                                                                                                                                                                                                                                                                                                                            8          8   2       v   2    e��     �   7   9   G      '            " X=" & to_string(x))) &LF&5��    7                 	   ~             	       5�_�                 8        ����                                                                                                                                                                                                                                                                                                                            8          8   2       v   2    e��     �   7   9   G      &            " X=" & to_string(x)) &LF&5��    7                      �                     5�_�                 8        ����                                                                                                                                                                                                                                                                                                                            8          8   2       v   2    e��   7 �   7   9   G      %            " X=" & to_string(x) &LF&5��    7                      �                     5�_�                 8       ����                                                                                                                                                                                                                                                                                                                            8          8   2       v   2    e�~     �   7   9   G      +            " X=" & character'image(x) &LF&5��    7          	          ~      	              �    7                     �                     �    7                                          �    7                 	   ~             	       �    7          	          ~      	              �    7                    ~                    5�_�                 8       ����                                                                                                                                                                                                                                                                                                                            8          8   2       v   2    e��     �   7   9   G      (            " X=" & string'image(x) &LF&5��    7          	          ~      	              5�_�                 8       ����                                                                                                                                                                                                                                                                                                                            8          8   2       v   2    e��     �   7   9   G      '            " X=" & stringimage(x) &LF&5��    7                     �                     5�_�                   8       ����                                                                                                                                                                                                                                                                                                                            8          8   2       v   2    e��   8 �   7   9   G      "            " X=" & string(x) &LF&5��    7                     �                     5�_�               8       ����                                                                                                                                                                                                                                                                                                                            8          :                 e�J     �   7   ;   G      6            " X=" & 'image(to_integer(signed(x))) &LF&   @            " Y=" & bit_vector'image(to_integer(signed(y))) &LF&   @            " Z=" & bit_vector'image(to_integer(signed(z))) &LF&�   7   9   G      @            " X=" & bit_vector'image(to_integer(signed(x))) &LF&5��    7                     ~                     �    8                     �                     �    9                     �                     �    7                     ~                     �    7                 
   ~             
       �    7          
          ~      
              �    7                 
   ~             
       �    8                  
   �              
       �    9                  
                  
       5�_�                 8   %    ����                                                                                                                                                                                                                                                                                                                            8          :                 e�Q     �   7   9   G      6            " X=" & bit_vector'image((signed(x))) &LF&5��    7   %       
           �      
               5�_�                 8   %    ����                                                                                                                                                                                                                                                                                                                            8          :                 e�S     �   7   9   G      5            " X=" & bit_vector'image(signed(x))) &LF&5��    7   %                  �                     5�_�                 8   .    ����                                                                                                                                                                                                                                                                                                                            8          :                 e�T     �   7   9   G      4            " X=" & bit_vector'image(signed(x)) &LF&5��    7   .                  �                     5�_�        	         8       ����                                                                                                                                                                                                                                                                                                                            8          :                 e�i     �   7   9   G      0            " X=" & signed'image(signed(x)) &LF&5��    7          
          ~      
              5�_�    
        	   8   %    ����                                                                                                                                                                                                                                                                                                                            8          :                 e�]     �   7   9   G      .            " X=" & bit_vector'image((x)) &LF&5��    7   %                  �                     5�_�  	            
   8   %    ����                                                                                                                                                                                                                                                                                                                            8          :                 e�]     �   7   9   G      -            " X=" & bit_vector'image(x)) &LF&5��    7   %                  �                     5�_�  
                 8   '    ����                                                                                                                                                                                                                                                                                                                            8          :                 e�^     �   7   9   G      ,            " X=" & bit_vector'image(x) &LF&5��    7   '                  �                     5�_�                         ����                                                                                                                                                                                                                                                                                                                                      F           V   6    e�9s     �              5��                          "                      5�_�   �   �   �   �   �   3       ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��^     �   2   4        5��    2                      �      a               5�_�   �   �           �   5        ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��_    �   5   6   <    �   5   6   <      `            assert false report "x is " & integer'image(to_integer(unsigned(Xv))) severity note;5��    5                      �              a       5�_�   �               �   6   M    ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��h     �   5   7   =      _            assert false report "x is " & integer'image(to_integer(unsigned(X))) severity note;5��    5   M                  <                     5�_�   �   �   �   �   �          ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��9     �         =      7        port map (x => xa, y => y, z => z, q => saida);5��                         `                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��=    �         =      .    signal xa, y, z : bit_vector(31 downto 0);5��                         u                     5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��C     �   *   ,   =                  xa <= Xv;5��    *                     (                     5�_�   �               �   3   M    ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��H    �   2   4   =      `            assert false report "x is " & integer'image(to_integer(unsigned(Xa))) severity note;5��    2   M                 +                    5�_�   �   �       �   �          ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e���     �         =      -    signal X, y, z : bit_vector(31 downto 0);5��                        t                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e���     �         =      -    signal X, Y, z : bit_vector(31 downto 0);5��                        w                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e���     �         =      -    signal X, Y, Z : bit_vector(31 downto 0);5��                        z                    �                        z                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e���     �         =      6        port map (x => X, y => y, z => z, q => saida);5��                        _                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e���     �         =      6        port map (x => X, y => Y, z => z, q => saida);5��                        g                    5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e���     �         =      6        port map (x => X, y => Y, z => Z, q => saida);5��       '                 o                    5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e���     �   *   ,   =                  X <= Xv;5��    *                    %                    5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e���     �   -   /   =                  Y <= Yv;5��    -                    {                    5�_�   �   �           �   1       ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e���    �   0   2   =                  Z <= Zv;5��    0                    �                    5�_�   �               �   3   L    ����                                                                                                                                                                                                                                                                                                                            ,          -          V       e��    �   2   4   =      _            assert false report "x is " & integer'image(to_integer(unsigned(X))) severity note;5��    2   L                 '                    5�_�   r           t   s   (   *    ����                                                                                                                                                                                                                                                                                                                            (          '   *       V   +    e��x     �   '   /        �   &   (   -      	        g5��    '                            �               �    &          "          �      "              5�_�   h           j   i          ����                                                                                                                                                                                                                                                                                                                            0   )       0   )       V   )    e��f     �              5��                          Y                      5�_�   b           d   c          ����                                                                                                                                                                                                                                                                                                                            -   )       -   )       V   )    e���     �         0       5��                          �                     �                          �                     �                          �                     5�_�   ^           `   _   !   $    ����                                                                                                                                                                                                                                                                                                                            +   )       +   )       V   )    e��Z     �       "   /      <        assert false report "BOT" & 'image(x) severity note;5��        $       
           @      
               5�_�   E   G       H   F          ����                                                                                                                                                                                                                                                                                                                               	                  V   	    e�ޯ     �      	        5��                          V       :               5�_�   F               G           ����                                                                                                                                                                                                                                                                                                                               	                  V   	    e�ޱ     �              5��                          V                      5�_�   5   7       8   6          ����                                                                                                                                                                                                                                                                                                                                                V       e��V     �         D      &    signal q: bit_vector(31 downto 0);5��                         �                      5�_�   6               7          ����                                                                                                                                                                                                                                                                                                                                                V       e��X     �   
      D      ,    signal x, y, z: bit_vector(31 downto 0);5��    
                     �                      5�_�   #           %   $   9       ����                                                                                                                                                                                                                                                                                                                            .   &       7          V   4    e�S,     �   8   :   O      	    end ;5��    8                     �                     5�_�                   '       ����                                                                                                                                                                                                                                                                                                                            N          N           V       e�Pc     �   '   (   K    �   &   (   K      9      file tb_file : text open read_mode is "alu_tb.dat";     variable tb_line: line;     variable space: character;   0  variable Av, Bv, res: bit_vector(63 downto 0);   : process is5��    &                     �                     �    &                     �              �       5�_�                           ����                                                                                                                                                                                                                                                                                                                            J          J           V       e�P8     �         K      use td.textio.all;5��                                               5�_�              	         .    ����                                                                                                                                                                                                                                                                                                                                                       e�Q     �         K      ?        (x"12345678", x"87654321", x"13579BDF",  -- Test case 55��       .                  �                     5��