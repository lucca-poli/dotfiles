Vim�UnDo� ��B�����șo�$'�A�d��L���xR�U                                      fں    _�                             ����                                                                                                                                                                                                                                                                                                                                                  V        fڹ    �                 library IEEE;   use IEEE.NUMERIC_BIT.all;       entity slow_clk is   
    port (           clk_in: in bit;           clk_out: out bit       );   end entity slow_clk;       architecture rtl of slow_clk is       )    signal counter: unsigned(9 downto 0);   (    signal current_state: bit := clk_in;          begin              timing: process(clk_in)   	    begin   #        if rising_edge(clk_in) then   #            counter <= counter + 1;   *            if counter = "1111111111" then   -                clk_out <= not current_state;               end if;           end if;       end process timing;          end architecture rtl;5��                                  7             5�_�                             ����                                                                                                                                                                                                                                                                                                                                                             fڰ     �               5��                                   (               5��