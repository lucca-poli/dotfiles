Vim�UnDo� ��Pp	\����g`������ׄ�C~��K  k   /    get_hout: adder32 port map (hv, hv, haso7);  5   !  �  �      �  �  �    fB�   � _�      �          �   �       ����                                                                                                                                                                                                                                                                                                                F                                      f4.     �   �   �  +    �   �   �  +    5��    �                      ]              D       5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                F           �          �          V       f4<     �   �   �  ,      C    signal av, bv, cv, dv, ev, fv, gv, hv: bit_vector(31 downto 0);5��    �                    i                    �    �                    p                    �    �                    w                    �    �   !                 ~                    �    �   (                 �                    �    �   /                 �                    �    �   6                 �                    �    �   =                 �                    �    �   G                 �                    5�_�  �  �          �   �   G    ����                                                                                                                                                                                                                                                                                                                F           �          �          V       f4D     �   �   �  ,      ^    signal a_out, b_out, c_out, d_out, e_out, f_out, g_out, h_out: bit__outector(31 downto 0);5��    �   G                  �                     5�_�  �  �          �   �   G    ����                                                                                                                                                                                                                                                                                                                F           �          �          V       f4D     �   �   �  ,      ]    signal a_out, b_out, c_out, d_out, e_out, f_out, g_out, h_out: bit_outector(31 downto 0);5��    �   G                  �                     5�_�  �  �          �   �   G    ����                                                                                                                                                                                                                                                                                                                F           �          �          V       f4E     �   �   �  ,      \    signal a_out, b_out, c_out, d_out, e_out, f_out, g_out, h_out: bit_utector(31 downto 0);5��    �   G                  �                     5�_�  �  �          �   �   G    ����                                                                                                                                                                                                                                                                                                                F           �          �          V       f4H     �   �   �  ,      [    signal a_out, b_out, c_out, d_out, e_out, f_out, g_out, h_out: bit_tector(31 downto 0);5��    �   G                  �                     5�_�  �  �          �   �   H    ����                                                                                                                                                                                                                                                                                                                F           �          �          V       f4I     �   �   �  ,      \    signal a_out, b_out, c_out, d_out, e_out, f_out, g_out, h_out: bit_vtector(31 downto 0);5��    �   H                  �                     5�_�  �  �          �   �   ,    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f4X     �   �   �  ,      .    get_aout: somador port map (h0, a_reg, a);�   �    ,      /    get_aout: somador port map (h0, a_reg, av);   /    get_bout: somador port map (h1, b_reg, bv);   /    get_cout: somador port map (h2, c_reg, cv);   /    get_dout: somador port map (h3, d_reg, dv);   /    get_eout: somador port map (h4, e_reg, ev);   /    get_fout: somador port map (h5, f_reg, fv);   /    get_gout: somador port map (h6, g_reg, gv);   /    get_hout: somador port map (hv, h_reg, hv);5��    �   ,                  9                     �    �   ,                  h                     �    �   ,                  �                     �    �   ,                  �                     �    �   ,                  �                     �    �   ,                  $                     �    �   ,                  S                     �    �   ,                  �                     �    �   ,                  9                     �    �   ,                  l                     �    �   ,                  �                     �    �   ,                  �                     �    �   ,                                       �    �   ,                  8                     �    �   ,                  k                     �    �   ,                  �                     5�_�  �  �          �  &       ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f4`     �  %  '  -                      �  %  '  ,    5��    %                     E!                     �    %                    E!                    �    %                    ]!                     5�_�  �  �          �  &       ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f4e     �  %  '  -                      done <= 5��    %                    ]!                     5�_�  �  �          �  &       ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f4e     �  %  '  -                      done <= ''5��    %                    ^!                     5�_�  �  �          �  &       ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f4g     �  &  (  .                      haso�  %  (  -                      done <= '1'5��    %                    `!                     �    %                   a!                     �    &                    r!                     �    &                    t!                     �    &                    s!                     �    &                   r!                    �    &                   r!                    �    &                	   r!             	       �    &                    z!                     5�_�  �  �          �  '       ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5b     �  &  (  .                      haso <= 5��    &                    y!                     �    &                   x!                    �    &                    {!                     �    &                    z!                     5�_�  �  �  �      �  '       ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5�     �  &  (  .                      haso <= 5��    &                     b!                     5�_�  �  �          �  '        ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5�     �  '  )  .    �  '  (  .    5��    '                     c!                     5�_�  �  �          �  (       ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5�     �  '  (                          haso <= 5��    '                     c!                     5�_�  �  �          �  '        ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5�     �  '  0  .    �  '  (  .    5��    '                     c!              �      5�_�  �  �          �  '        ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5�     �  &  '           5��    &                     b!                     5�_�  �  �          �  '        ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5�     �  &  (  5      Z        inst6: somador port map (a => aout, b => x"6a09e667",  soma => haso(31 downto 0));5��    &          3           b!      3               5�_�  �  �          �  '        ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5�     �  &  (  5      '6a09e667",  soma => haso(31 downto 0));5��    &          	           b!      	               5�_�  �  �          �  '        ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5�     �  &  (  5      ,  soma => haso(31 downto 0));5��    &                     b!                     5�_�  �  �          �  '        ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5�     �  &  (  5      haso(31 downto 0));5��    &                     b!                     5�_�  �  �          �  '   #    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5�     �  &  (  5      #                haso(31 downto 0));5��    &  "                  �!                     �    &  !              	   �!             	       5�_�  �  �          �  (        ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5�     �  '  )  5      [        inst7: somador port map (a => bout, b => x"bb67ae85",  soma => haso(63 downto 32));5��    '          G          �!      G              �    '  "              	   �!             	       5�_�  �  �          �  )        ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5�     �  -  /  5      ^        inst13: somador port map (a => hout, b => x"5be0cd19",  soma => haso(255 downto 224));�  ,  .  5      ^        inst12: somador port map (a => gout, b => x"1f83d9ab",  soma => haso(223 downto 192));�  +  -  5      ^        inst11: somador port map (a => fout, b => x"9b05688c",  soma => haso(191 downto 160));�  *  ,  5      ^        inst10: somador port map (a => eout, b => x"510e527f",  soma => haso(159 downto 128));�  )  +  5      \        inst9: somador port map (a => dout, b => x"a54ff53a",  soma => haso(127 downto 96));�  (  *  5      [        inst8: somador port map (a => cout, b => x"3c6ef372",  soma => haso(95 downto 64));5��    (          G          �!      G              �    (  "              	   �!             	       �    )          G          �!      G              �    )  #              	   "             	       �    *          H          "      H              �    *  $              	   6"             	       �    +          H          @"      H              �    +  $              	   d"             	       �    ,          H          n"      H              �    ,  $              	   �"             	       �    -          H          �"      H              �    -  $              	   �"             	       5�_�  �  �          �  '   %    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5�     �  &  (  5      *                haso(31 downto 0) <= _out;5��    &  %                  �!                     5�_�  �  �          �  '   "    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6     �  &  (  5      +                haso(31 downto 0) <= a_out;5��    &  "                  �!                     5�_�  �  �          �  (   #    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6     �  '  )  5      +                haso(63 downto 32) <= _out;5��    '  #                  �!                     5�_�  �  �          �  )   #    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6     �  (  *  5      +                haso(95 downto 64) <= _out;5��    (  #                  �!                     5�_�  �  �          �  *   $    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6     �  )  +  5      ,                haso(127 downto 96) <= _out;5��    )  $                  "                     5�_�  �  �          �  (   (    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6
     �  '  )  5      -                haso(63 downto 32)   <= _out;5��    '  (                  �!                     5�_�  �  �          �  )   (    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6     �  (  *  5      -                haso(95 downto 64)   <= _out;5��    (  (                  �!                     5�_�  �  �          �  *   (    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6     �  )  +  5      -                haso(127 downto 96)  <= _out;5��    )  (                  "                     5�_�  �  �          �  +   (    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6     �  *  ,  5      -                haso(159 downto 128) <= _out;5��    *  (                  F"                     5�_�  �  �          �  ,   (    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6     �  +  -  5      -                haso(191 downto 160) <= _out;5��    +  (                  u"                     5�_�  �  �          �  -   (    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6     �  ,  .  5      -                haso(223 downto 192) <= _out;5��    ,  (                  �"                     5�_�  �  �          �  .   (    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6     �  -  /  5      -                haso(255 downto 224) <= _out;5��    -  (                  �"                     5�_�  �  �          �  %       ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6J     �  $  &  5      %            elsif iteration = 63 then5��    $                    1!                     5�_�  �  �  �      �  %       ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6g   ? �  $  &  5      &            elsif (iteration = 63 then5��    $                    1!                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f7^   A �        5      %        q: out bit_vector(7 downto 0)5��                        v                     5�_�  �  �          �   O       ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f7�   C �   N   P  5      )            q: out bit_vector(7 downto 0)5��    N                    �                    5�_�  �  �          �   6       ����                                                                                                                                                                                                                                                                                                                F           �          �   %       V   9    f<     �   9   ;  9      use IEEE.numeric_std.all;�   7   ;  7      ieee�   6   9  6       �   6   8  5    5��    6                      q                     �    6                      q                     �    7                      r                     �    7                     t                     �    7                     s                     �    7                     r                    �    7                     r                    �    7                     r                    �    7                      r                     �    7                     r              D       �    9                      �                      5�_�  �  �          �   6       ����                                                                                                                                                                                                                                                                                                                J           �          �   %       V   9    f<     �   6   8  :       �   6   8  9    5��    6                      q                     �    6                      q                     �    6                     q                    �    6                     q                    �    6   
                  {                     �    6   	                 z                    �    6   
                  {                     �    6   	                 z                    �    6                     |                     �    6   
                  {                     �    6   	                 z                    �    6                     �                     �    6                     �                     �    6                     �                     �    6                     �                     �    6                     �                     �    6                                          �    6                     ~                     �    6                     }                     �    6                     |                     �    6   
                  {                     �    6   	                 z                    �    6                     �                     �    6                     �                     �    6                     �                     �    6                     �                     �    6                     �                     �    6                     �                     �    6                     �                     �    6                     �                     �    6                     �                     �    6                     �                     �    6                                          �    6                     ~                     �    6                     }                     �    6                     |                     �    6   
                  {                     �    6   	                 z                    �    6   	                 z                    �    6   	                 z                    5�_�  �  �          �   7       ����                                                                                                                                                                                                                                                                                                                K           �          �   %       V   9    f<1     �   6   8  :      use IEEE.IEEE_BIT_CONTEXT5��    6                     �                     �    6                    �                    5�_�  �  �          �   7       ����                                                                                                                                                                                                                                                                                                                K           �          �   %       V   9    f<8     �   6   7          use IEEE.IEEE_BIT_CONTEXT.ALL;5��    6                      q                     5�_�  �  �          �   8        ����                                                                                                                                                                                                                                                                                                                J           �          �   %       V   9    f<:   F �   7   8          library IEEE;   use IEEE.std_logic_1164.all;   use IEEE.numeric_std.all;    5��    7                      r      F               5�_�  �  �  �      �          ����                                                                                                                                                                                                                                                                                                                F                     5           V        f=�     �        5    5��                          �                     5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                G                     6           V        f=�   G �      +  6    �        6    5��                          �                    5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                Z                     +           V       f>#   I �                entity somador is   
    port (   '        A : in bit_vector(31 downto 0);   '        B : in bit_vector(31 downto 0);   '        S : out bit_vector(31 downto 0)       );   end entity somador;       %architecture behavioral of somador is   +    signal carry : bit_vector(31 downto 0);   begin   "    sum: for i in 0 to 30 generate   +        S(i) <= A(i) xor B(i) xor carry(i);   T        carry(i+1) <= (A(i) and B(i)) or (A(i) and carry(i)) or (B(i) and carry(i));       end generate;       +    S(31) <= A(31) xor B(31) xor carry(31);          end architecture behavioral;    5��                          �                    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                F                                    f@�   K �      5          a <= h0;�      5          a_reg <= h0;       b_reg <= h1;       c_reg <= h2;       d_reg <= h3;       e_reg <= h4;       f_reg <= h5;       g_reg <= h6;       h_reg <= h7;5��                        %                      �                        2                      �                        ?                      �                        L                      �                        Y                      �                        f                      �                        s                      �                        �                      �                        %                      �                        3                      �                        A                      �                        O                      �                        ]                      �                        k                      �                        y                      �                        �                      5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                F                                    fAj     �   �   �  5    �   �   �  5    5��    �                      _              \       5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                F                                    fAr     �   �   �  6      [    signal a_reg, b_reg, c_reg, d_reg, e_reg, f_reg, g_reg, h_reg: bit_vector(31 downto 0);5��    �          1                 1               5�_�  �  �          �   �   )    ����                                                                                                                                                                                                                                                                                                                F                                    fAx     �   �   �  6      *    signal a_reg: bit_vector(31 downto 0);5��    �   )                  ,                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                F                                    fA�     �   �   �  6      [    signal a_reg, b_reg, c_reg, d_reg, e_reg, f_reg, g_reg, h_reg: bit_vector(31 downto 0);5��    �                     ?                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                F                                    fA�     �   �   �  6      V    signal , b_reg, c_reg, d_reg, e_reg, f_reg, g_reg, h_reg: bit_vector(31 downto 0);5��    �                     ?                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                F                                    fA�     �   �   �          T    signal b_reg, c_reg, d_reg, e_reg, f_reg, g_reg, h_reg: bit_vector(31 downto 0);5��    �                      4      U               5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                F                                    fA�     �   �   �  5    �   �   �  5    5��    �                      4              1       5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                F                                    fA�     �   �   �  6    �   �   �  6    5��    �                      e              1       5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                F                                    fA�     �   �   �  7    �   �   �  7    5��    �                      �              1       5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                F                                     fA�     �   �   �  8    �   �   �  8    5��    �                      �              1       5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                F                   !                 fA�     �   �   �  9    �   �   �  9    5��    �                      �              1       5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                F                   "                 fA�     �   �   �  :    �   �   �  :    5��    �                      )              1       5�_�  �             �   �       ����                                                                                                                                                                                                                                                                                                                F                   #                 fA�     �   �   �  ;    �   �   �  ;    5��    �                      Z              1       5�_�  �                �       ����                                                                                                                                                                                                                                                                                                                F                   $                 fA�     �   �   �  <    �   �   �  <    5��    �                      �              1       5�_�                  �       ����                                                                                                                                                                                                                                                                                                                F                   %                 fA�     �   �   �  =      0    signal a_reg: bit_vector(31 downto 0) := h0;5��    �                    ?                    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                F                   %                 fA�     �   �   �  =      0    signal a_reg: bit_vector(31 downto 0) := h0;5��    �                    p                    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                F                   %                 fA�     �   �   �  =      0    signal a_reg: bit_vector(31 downto 0) := h0;5��    �                    �                    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                F                   %                 fA�     �   �   �  =      0    signal a_reg: bit_vector(31 downto 0) := h0;5��    �                    �                    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                F                   %                 fA�     �   �   �  =      0    signal a_reg: bit_vector(31 downto 0) := h0;5��    �                                        5�_�                 �       ����                                                                                                                                                                                                                                                                                                                F                   %                 fA�     �   �   �  =      0    signal a_reg: bit_vector(31 downto 0) := h0;5��    �                    4                    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                F                   %                 fA�     �   �   �  =      0    signal a_reg: bit_vector(31 downto 0) := h0;5��    �                    e                    5�_�    	             �       ����                                                                                                                                                                                                                                                                                                                F                   %                 fA�     �   �   �          0    signal a_reg: bit_vector(31 downto 0) := h0;5��    �                      �      1               5�_�    
          	   �   .    ����                                                                                                                                                                                                                                                                                                                F           �   .       �   .          .    fA�   L �   �   �  <      0    signal b_reg: bit_vector(31 downto 0) := h0;   0    signal c_reg: bit_vector(31 downto 0) := h0;   0    signal d_reg: bit_vector(31 downto 0) := h0;   0    signal e_reg: bit_vector(31 downto 0) := h0;   0    signal f_reg: bit_vector(31 downto 0) := h0;   0    signal g_reg: bit_vector(31 downto 0) := h0;   0    signal h_reg: bit_vector(31 downto 0) := h0;5��    �   .                 b                    �    �   .                 �                    �    �   .                 �                    �    �   .                 �                    �    �   .                 &                    �    �   .                 W                    �    �   .                 �                    5�_�  	            
          ����                                                                                                                                                                                                                                                                                                                F           �   .       �   .          .    fA�   M �           	       av <= h0;       bv <= h1;       cv <= h2;       dv <= h3;       ev <= h4;       fv <= h5;       gv <= h6;       hv <= h7;    5��          	               L!      q               5�_�  
                      ����                                                                                                                                                                                                                                                                                                                F           �   .       �   .          .    fG�     �         3    5��                                                  5�_�                         ����                                                                                                                                                                                                                                                                                                                G           �   .       �   .          .    fG�     �        7      use IEEE.numeric_std.all;�         5       �         4    5��                                                  �                                                  �                                                �                                                �                                                �                                                �                                                �                                                  �                                          D       �                          D                       5�_�                        ����                                                                                                                                                                                                                                                                                                                J           �   .       �   .          .    fG�     �                use IEEE.std_logic_1164.all;5��                                                5�_�                    	    ����                                                                                                                                                                                                                                                                                                                I           �   .       �   .          .    fG�   N �        6      use IEEE.numeric_std.all;5��       	                                      �                                               �                                               �                                               �       
                                        �       	                                      �                                               �                                               �       
                                        �       	                                      �       	                                      �       	                                      5�_�                 ^        ����                                                                                                                                                                                                                                                                                                                I                                V       fH�     �  	            2    get_hout: somador port map (hv, h_reg, h_out);�    
          2    get_gout: somador port map (h6, g_reg, g_out);�    	          2    get_fout: somador port map (h5, f_reg, f_out);�              2    get_eout: somador port map (h4, e_reg, e_out);�              2    get_dout: somador port map (h3, d_reg, d_out);�              2    get_cout: somador port map (h2, c_reg, c_out);�              2    get_bout: somador port map (h1, b_reg, b_out);�              2    get_aout: somador port map (h0, a_reg, a_out);�   �   �          0        	make1: somador port map(op1, op2, op3);�   �   �          8        	make5: somador port map(op4, w_vec(i-16), op5);�   �   �          0        	make4: somador port map(op3, op2, op4);�   �   �          7        	make3: somador port map(op3, w_vec(i-7), op3);�   ]   _  6          component somador  is5��    ]                    d                    �    �                    �                    �    �                    �                    �    �                                        �    �                    $                    �                       r                    �                       �                    �                       �                    �                                           �                       >                    �                       q                    �                       �                    �    	                   �                    5�_�                 `       ����                                                                                                                                                                                                                                                                                                                I                                V       fH�     �   _   a  6      +            A : in bit_vector(31 downto 0);5��    _                    �                    5�_�                 a       ����                                                                                                                                                                                                                                                                                                                I                                V       fH�     �   `   b  6      +            B : in bit_vector(31 downto 0);5��    `                    �                    5�_�                 b       ����                                                                                                                                                                                                                                                                                                                I                                V       fH�   O �   a   c  6      +            S : out bit_vector(31 downto 0)5��    a                    �                    5�_�                 !   
    ����                                                                                                                                                                                                                                                                                                                I                                V       fJ�     �       !          =        rst : in bit;                          -- Reset input5��                           `      >               5�_�                         ����                                                                                                                                                                                                                                                                                                                H                                V       fJ�     �      !  5      ?        clk : in bit;                            -- Clock input5��                         +                     �                         7                     �                         6                     �                        5                    5�_�                 ,       ����                                                                                                                                                                                                                                                                                                                H                                V       fJ�     �   +   -  6              �   +   -  5    5��    +                      N              	       �    +                     V                     5�_�                 ,       ����                                                                                                                                                                                                                                                                                                                I                                V       fJ�     �   +   -  6              if enable = 5��    +                     b                     5�_�                 ,       ����                                                                                                                                                                                                                                                                                                                I                                V       fJ�     �   +   -  6              if enable = ''5��    +                     c                     5�_�                 ,       ����                                                                                                                                                                                                                                                                                                                I                                V       fJ�     �   +   -  6              if enable = '1'5��    +                     e                     �    +                    f                    5�_�                 -       ����                                                                                                                                                                                                                                                                                                                I           -          1                 fJ�     �   -   2  6      '            counter <= (others => '0');   #        elsif rising_edge(clk) then   #            counter <= counter + 1;           end if;�   ,   .  6              if rst = '1' then5��    ,                     s                     �    -                     �                     �    .                     �                     �    /                     �                     �    0                                          5�_�                 1       ����                                                                                                                                                                                                                                                                                                                I           -          1                 fJ�     �   1   3  7                  �   1   3  6    5��    1                                           �    1                     %                     �    1                    '                    �    1                                         �    1                     %                     �    1                    '                    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fK&     �   �   �  8          �   �   �  7    5��    �                      �                     �    �                     �                     �    �                                        5�_�                 �       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fK=     �   �   �  8          signal done: bit := 0;5��    �                                          5�_�                 �       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fK=     �   �   �  8          signal done: bit := ;5��    �                                          5�_�                 �       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fK>     �   �   �  8          signal done: bit := '';5��    �                                          5�_�                  �       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fKC     �   �   �  8          signal done: bit := '0';5��    �                                        5�_�    !              �   -    ����                                                                                                                                                                                                                                                                                                                J           -          1                 fKT   P �   �   �  8      9    counter: counter_6bit port map (clk, rst, iteration);5��    �   -                  �                     �    �   .                 �                    �    �   .                 �                    �    �   .                 �                    5�_�     "          !   Z       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fK�     �   Y   Z          A            rst : in bit;                          -- Reset input5��    Y                      �      B               5�_�  !  #          "   Y       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fK�   Q �   X   Z  7      C            clk : in bit;                            -- Clock input5��    X                     �                     �    X                    �                    �    X                    �                    5�_�  "  $          #  &       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fK�     �  &  (  8                      �  &  (  7    5��    &                     �!                     �    &                    �!                     �    &                    "                     �    &                     "                     �    &                   �!                    �    &                   �!                    �    &                
   �!             
       5�_�  #  %          $  '       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fK�     �  &  (  8                      enable <= 5��    &                    	"                     5�_�  $  &          %  '       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fK�     �  &  (  8                      enable <= ''5��    &                    
"                     5�_�  %  '          &  '       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fK�     �  &  (  8                      enable <= '0'5��    &                    "                     5�_�  &  (          '  )       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fK�     �  )  +  9                      �  )  +  8    5��    )                     Q"                     �    )                    a"                     �    )                    c"                     �    )                    b"                     �    )                   a"                    �    )                   a"                    �    )                
   a"             
       5�_�  '  )          (  *       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fK�     �  )  +  9                      enable <= 5��    )                    k"                     5�_�  (  *          )  *       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fK�     �  )  +  9                      enable <= ''5��    )                    l"                     5�_�  )  +          *  *       ����                                                                                                                                                                                                                                                                                                                J           -          1                 fK�   R �  )  +  9                      enable <= '1'5��    )                    n"                     5�_�  *  ,          +  3       ����                                                                                                                                                                                                                                                                                                                J                             v       fL     �  4  6  ;                  current_kpw�  3  6  :                  �  3  5  9    5��    3                     �#                     �    3                     �#                     �    3                    �#                     �    4                    	$                     �    4                    $                     �    4                    $                     �    4                    
$                     �    4                   	$                    �    4                   	$                    �    4                   	$                    �    4                    $                     �    4                   $                    �    4                    $                     �    4                    $                     �    4                   $                    �    4  !                  $                     �    4                     $                     �    4                    $                     �    4                    $                     �    4                    $                     �    4                    $                     �    4                   $                    �    4                   $                    �    4                   $                    5�_�  +  -          ,  5   "    ����                                                                                                                                                                                                                                                                                                                J                             v       fL%     �  4  6  ;      "            current_kpw <= kpw_vec5��    4  "                  $                     5�_�  ,  .          -  5   #    ����                                                                                                                                                                                                                                                                                                                J                             v       fL&     �  4  6  ;      $            current_kpw <= kpw_vec()5��    4  #                   $                     �    4  #              	    $             	       �    4  #       	           $      	              �    4  #              	    $             	       5�_�  -  /          .  5   -    ����                                                                                                                                                                                                                                                                                                                J                             v       fL(   S �  4  6  ;      -            current_kpw <= kpw_vec(iteration)5��    4  -                  *$                     5�_�  .  0          /  '       ����                                                                                                                                                                                                                                                                                                                J                             v       fL�     �  &  '                          enable <= '0';5��    &                     �!                     5�_�  /  1          0  )       ����                                                                                                                                                                                                                                                                                                                J                             v       fL�     �  (  )                          enable <= '1';5��    (                     2"                     5�_�  0  2          1           ����                                                                                                                                                                                                                                                                                                                J                             v       fL�     �      !  9      L        clk, rst, enable : in bit;                            -- Clock input5��                         2                     5�_�  1  3          2           ����                                                                                                                                                                                                                                                                                                                J                             v       fL�     �      !  9      E        clk, rst, : in bit;                            -- Clock input5��                         0                     5�_�  2  4          3   ,       ����                                                                                                                                                                                                                                                                                                                J                             v       fL�     �   +   ,                  if enable = '1' then5��    +                      E                     5�_�  3  5          4   1       ����                                                                                                                                                                                                                                                                                                                I                             v       fL�     �   0   1                  end if;5��    0                      �                     5�_�  4  6          5   ,       ����                                                                                                                                                                                                                                                                                                                H           0          ,                 fL�     �   +   -  7                  if rst = '1' then5��    +                     M                     5�_�  5  7          6   -       ����                                                                                                                                                                                                                                                                                                                H           0          ,                 fL�     �   ,   .  7      +                counter <= (others => '0');5��    ,                     k                     5�_�  6  8          7   .       ����                                                                                                                                                                                                                                                                                                                H           0          ,                 fL�     �   -   /  7      '            elsif rising_edge(clk) then5��    -                     �                     5�_�  7  9          8   /       ����                                                                                                                                                                                                                                                                                                                H           0          ,                 fL�     �   .   0  7      '                counter <= counter + 1;5��    .                     �                     5�_�  8  :          9   0       ����                                                                                                                                                                                                                                                                                                                H           0          ,                 fL�     �   /   1  7                  end if;5��    /                     �                     5�_�  9  ;          :   W       ����                                                                                                                                                                                                                                                                                                                H           0          ,                 fL�     �   V   X  7      P            clk, rst, enable : in bit;                            -- Clock input5��    V                     F                     5�_�  :  <          ;   W       ����                                                                                                                                                                                                                                                                                                                H           0          ,                 fL�     �   V   X  7      I            clk, rst, : in bit;                            -- Clock input5��    V                     D                     5�_�  ;  =          <   �       ����                                                                                                                                                                                                                                                                                                                H           0          ,                 fL�     �   �   �              signal enable: bit := '0';5��    �                      p                     5�_�  <  >          =   �   .    ����                                                                                                                                                                                                                                                                                                                H           0          ,                 fL�   U �   �   �  6      A    counter: counter_6bit port map (clk, rst, enable, iteration);5��    �   .                  .                     5�_�  =  ?          >   �        ����                                                                                                                                                                                                                                                                                                                H           �   /       �   0       V   V    fM     �   �   �  6    �   �   �  6    5��    �                      �              �      5�_�  >  @          ?   �       ����                                                                                                                                                                                                                                                                                                                H           �          �                 fM     �   �   �  >      ,    signal a: bit_vector(31 downto 0) := h0;�   �   �  >      0    signal a_reg: bit_vector(31 downto 0) := h0;   0    signal b_reg: bit_vector(31 downto 0) := h1;   0    signal c_reg: bit_vector(31 downto 0) := h2;   0    signal d_reg: bit_vector(31 downto 0) := h3;   0    signal e_reg: bit_vector(31 downto 0) := h4;   0    signal f_reg: bit_vector(31 downto 0) := h5;   0    signal g_reg: bit_vector(31 downto 0) := h6;   0    signal h_reg: bit_vector(31 downto 0) := h7;5��    �                     �                     �    �                     �                     �    �                                          �    �                     G                     �    �                     t                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                                          �    �                     J                     �    �                     x                     �    �                     �                     �    �                     �                     �    �                                          5�_�  ?  A          @   �       ����                                                                                                                                                                                                                                                                                                                H           �          �                 fM   V �   �   �          C    signal av, bv, cv, dv, ev, fv, gv, hv: bit_vector(31 downto 0);5��    �                      p      D               5�_�  @  B          A     +    ����                                                                                                                                                                                                                                                                                                                H             +         /          /    fYg     �      =   	   -    get_aout: adder32 port map (h0, a_reg, );   -    get_bout: adder32 port map (h1, b_reg, );   -    get_cout: adder32 port map (h2, c_reg, );   -    get_dout: adder32 port map (h3, d_reg, );   -    get_eout: adder32 port map (h4, e_reg, );   -    get_fout: adder32 port map (h5, f_reg, );   -    get_gout: adder32 port map (h6, g_reg, );   -    get_hout: adder32 port map (hv, h_reg, );    �    	  =    �      =      2    get_aout: adder32 port map (h0, a_reg, a_out);   2    get_bout: adder32 port map (h1, b_reg, b_out);   2    get_cout: adder32 port map (h2, c_reg, c_out);   2    get_dout: adder32 port map (h3, d_reg, d_out);   2    get_eout: adder32 port map (h4, e_reg, e_out);   2    get_fout: adder32 port map (h5, f_reg, f_out);   2    get_gout: adder32 port map (h6, g_reg, g_out);   2    get_hout: adder32 port map (hv, h_reg, h_out);5��      +                  C                     �      +                  q                     �    	  +                  �                     �    
  +                  �                     �      +                  �                     �      +                  )                      �      +                  W                      �      +                  �                      �      +                  C                     �      +                  �                     �    	  +                  �                     �    
  +                                        �      +                  S                      �      +                  �                      �      +                  �                      �      +                  !                     5�_�  A  C          B  -        ����                                                                                                                                                                                                                                                                                                                H          -   +      4   +       V   +    fY|     �  ,  -          .                haso(31 downto 0)    <= a_out;   .                haso(63 downto 32)   <= b_out;   .                haso(95 downto 64)   <= c_out;   .                haso(127 downto 96)  <= d_out;   .                haso(159 downto 128) <= e_out;   .                haso(191 downto 160) <= f_out;   .                haso(223 downto 192) <= g_out;   .                haso(255 downto 224) <= h_out;5��    ,                     l#      x              5�_�  B  D          C     <    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �    	  5      C    get_aout: adder32 port map (h0, a_reg, haso(31 downto 0));   );5��      <                  T                     5�_�  C  E          D     <    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �    	  5      B    get_aout: adder32 port map (h0, a_reg, haso(31 downto 0);   );5��      <                  T                     5�_�  D  F          E     <    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �    	  5      A    get_aout: adder32 port map (h0, a_reg, haso(31 downto 0)   );5��      <                  T                     5�_�  E  G          F  	   =    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �    
  5      C    get_bout: adder32 port map (h1, b_reg, haso(63 downto 32));  );5��      =                  �                     5�_�  F  H          G  	   =    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �    
  5      B    get_bout: adder32 port map (h1, b_reg, haso(63 downto 32);  );5��      =                  �                     5�_�  G  I          H  	   =    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �    
  5      A    get_bout: adder32 port map (h1, b_reg, haso(63 downto 32)  );5��      =                  �                     5�_�  H  J          I  
   =    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �  	    5      C    get_cout: adder32 port map (h2, c_reg, haso(95 downto 64));  );5��    	  =                  �                     5�_�  I  K          J  
   =    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �  	    5      B    get_cout: adder32 port map (h2, c_reg, haso(95 downto 64);  );5��    	  =                  �                     5�_�  J  L          K  
   =    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �  	    5      A    get_cout: adder32 port map (h2, c_reg, haso(95 downto 64)  );5��    	  =                  �                     5�_�  K  M          L     >    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �  
    5      C    get_dout: adder32 port map (h3, d_reg, haso(127 downto 96)); );5��    
  >                                        5�_�  L  N          M     >    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �  
    5      B    get_dout: adder32 port map (h3, d_reg, haso(127 downto 96); );5��    
  >                                        5�_�  M  O          N     >    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �  
    5      A    get_dout: adder32 port map (h3, d_reg, haso(127 downto 96) );5��    
  >                                        5�_�  N  P          O     ?    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �      5      C    get_eout: adder32 port map (h4, e_reg, haso(159 downto 128)););5��      ?                  W                      5�_�  O  Q          P     ?    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �      5      B    get_eout: adder32 port map (h4, e_reg, haso(159 downto 128););5��      ?                  W                      5�_�  P  R          Q     ?    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �      5      C    get_fout: adder32 port map (h5, f_reg, haso(191 downto 160)););5��      ?                  �                      5�_�  Q  S          R     ?    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �      5      B    get_fout: adder32 port map (h5, f_reg, haso(191 downto 160););5��      ?                  �                      5�_�  R  T          S     ?    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �      5      C    get_gout: adder32 port map (h6, g_reg, haso(223 downto 192)););5��      ?                  �                      5�_�  S  U          T     ?    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �      5      B    get_gout: adder32 port map (h6, g_reg, haso(223 downto 192););5��      ?                  �                      5�_�  T  V          U     ?    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�     �      5      C    get_hout: adder32 port map (hv, h_reg, haso(255 downto 224)););5��      ?                  !                     5�_�  U  W          V     ?    ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�   W �      5      B    get_hout: adder32 port map (hv, h_reg, haso(255 downto 224););5��      ?                  !                     5�_�  V  �          W   �       ����                                                                                                                                                                                                                                                                                                                H          -   +      -   +       V   +    fY�   g �   �   �          [    signal a_out, b_out, c_out, d_out, e_out, f_out, g_out, h_out: bit_vector(31 downto 0);5��    �                      h      \               5�_�  W  �  X      �  4        ����                                                                                                                                                                                                                                                                                                                H           �          �                 f��     �  4            �  4            5��    4                     z#              �      5�_�  �  �          �  5       ����                                                                                                                                                                                                                                                                                                                H           �          �                 f��     �  4  6  F      entity somador32 is5��    4         	          �#      	              5�_�  �  �          �  :       ����                                                                                                                                                                                                                                                                                                                H           �          �                 f��     �  9  ;  F      end somador32;5��    9         	          �#      	              5�_�  �  �          �  <       ����                                                                                                                                                                                                                                                                                                                H           �          �                 f��   h �  ;  =  F      'architecture behavioral of somador32 is5��    ;         	          $      	              5�_�  �  �          �   `       ����                                                                                                                                                                                                                                                                                                                H           �          �                 f�9   i �   _   a  F      +            r : out bit_vector(31 downto 0)5��    _                    k                    5�_�  �  �          �  $       ����                                                                                                                                                                                                                                                                                                                H                    F          V       f��     �  #  %  F          process(clk)5��    #                    L"                     5�_�  �  �          �  &        ����                                                                                                                                                                                                                                                                                                                H                    F          V       f��     �  %  '  F       5��    %                     ]"                     �    %                   j"                    5�_�  �  �          �  &       ����                                                                                                                                                                                                                                                                                                                H                    F          V       f��     �  %  '  F              if rst = 5��    %                    n"                     5�_�  �  �          �  &       ����                                                                                                                                                                                                                                                                                                                H                    F          V       f��     �  %  '  F              if rst = ''5��    %                    o"                     5�_�  �  �          �  &       ����                                                                                                                                                                                                                                                                                                                H                    F          V       f��     �  %  '  F              if rst = '1'5��    %                    q"                     �    %                   r"                    �    %                   r"                    �    %                   r"                    5�_�  �  �          �  '       ����                                                                                                                                                                                                                                                                                                                H                    F          V       f��     �  &  (  F               if rising_edge(clk) then5��    &                    "                     5�_�  �  �          �  &       ����                                                                                                                                                                                                                                                                                                                H                    F          V       f��     �  %  (  F              if rst = '1' then5��    %                   v"              	       �    &                    w"                    �    &                   �"                    5�_�  �  �          �  '       ����                                                                                                                                                                                                                                                                                                                H                    G          V       f��     �  &  (  G                  done <= 5��    &                    �"                     5�_�  �  �          �  '       ����                                                                                                                                                                                                                                                                                                                H                    G          V       f��     �  &  (  G                  done <= ''5��    &                    �"                     5�_�  �  �          �  '       ����                                                                                                                                                                                                                                                                                                                H                    G          V       f��     �  &  (  G                  done <= '0'5��    &                    �"                     5�_�  �  �          �  *       ����                                                                                                                                                                                                                                                                                                                H                    G          V       f��     �  (  *  G                  if rst = '1' then    �  )  +  G                      done <= '0';5��    )                    �"                     �    )                    �"                     �    )                    �"                     �    )                    �"                     �    )                    �"                     �    )                    �"                     �    )                    �"                     �    )                    �"                     �    )                    �"                     �    )                    �"                     �    )                    �"                     �    )                    �"                     �    )                    �"                     �    )                    �"                     �    )                    �"                     �    )                    �"                     �    )                    �"                     �    )  
                  �"                     �    )  	                  �"                     �    )          	           �"      	               �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                    �"                     �    (                   �"                    �    (                    �"                     �    (                    �"                     5�_�  �  �          �  )       ����                                                                                                                                                                                                                                                                                                                H                    F          V       f��     �  (  )                      5��    (                     �"                     5�_�  �  �  �      �  )       ����                                                                                                                                                                                                                                                                                                                H                    E          V       f��     �  (  *  E      %            elsif iteration = 63 then5��    (                   �"                    5�_�  �  �          �  )       ����                                                                                                                                                                                                                                                                                                                H                    E          V       f��   j �  (  *  E      %           ielsif iteration = 63 then5��    (                   �"                    �    (                    �"                    5�_�  �  �          �  '       ����                                                                                                                                                                                                                                                                                                                H                    E          V       f�     �  '  )  F                  �  '  )  E    5��    '                     �"                     �    '                    �"                     5�_�  �  �          �  (       ����                                                                                                                                                                                                                                                                                                                H                    F          V       f�     �  '  )  F                  iter5��    '                    �"                     5�_�  �  �          �  (       ����                                                                                                                                                                                                                                                                                                                H                    F          V       f�     �  '  )  F                  iter[]5��    '                    �"                     �    '                    �"                     �    '                    �"                     �    '                    �"                     �    '                    �"                     �    '                	   �"             	       �    '         	          �"      	              �    '                	   �"             	       5�_�  �  �          �  (       ����                                                                                                                                                                                                                                                                                                                H                    F          V       f�     �  '  )  F                  iteration5��    '                     �"                     5�_�  �  �          �  (        ����                                                                                                                                                                                                                                                                                                                H                    F          V       f�     �  '  (           5��    '                     �"                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                H                               V       f�     �        E    5��                          �                     5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                I                               V       f�     �      4  F    �        F    5��                          �              �      5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                b                               V       f�     �        _      entity reg32 is5��                     	                	       �                                            �                                            �                                            �              	                	              5�_�  �  �          �   !   %    ����                                                                                                                                                                                                                                                                                                                b                               V       f�2     �       "  `          �       "  _    5��                           :              	       �                          :                    �                          E                     �        
                 D                    �                          E                     �        
                  D                     �        	                  C                     �                         B                    �                      
   K             
       �               
          K      
              �                      
   K             
       5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                c                               V       f�K     �       "  `              data: in bit_vector5��                          U                     5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                c                               V       f�L     �       "  `              data: in bit_vector()5��                          V                     5�_�  �  �          �   !   (    ����                                                                                                                                                                                                                                                                                                                c                               V       f�P     �       "  `      (        data: in bit_vector(31 downto 0)5��        (                  b                     5�_�  �  �          �   "       ����                                                                                                                                                                                                                                                                                                                c                               V       f�S     �   !   #  `      &        d: in bit_vector(31 downto 0);5��    !                    }                    �    !                                        5�_�  �  �          �   #       ����                                                                                                                                                                                                                                                                                                                c                               V       f�[     �   "   $  `      &        q: out bit_vector(31 downto 0)5��    "                    �                    5�_�  �  �          �   %       ����                                                                                                                                                                                                                                                                                                                c                               V       f�_     �   $   &  `      end entity reg32;5��    $                    �                    �    $                     �                     �    $                     �                     �    $                    �                    �    $                    �                    �    $                    �                    5�_�  �  �          �   '       ����                                                                                                                                                                                                                                                                                                                c                               V       f�c     �   &   (  `      !architecture Behavior of reg32 is5��    &                    �                    �    &                     �                     �    &                     �                     �    &                    �                    �    &                    �                    �    &                    �                    5�_�  �  �          �   0       ����                                                                                                                                                                                                                                                                                                                c                               V       f�r     �   /   1  `                  Q <= D;5��    /                     �                     5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                c                               V       f��     �      !  `              rst, clk: in bit;5��                         0                     5�_�  �  �          �   0       ����                                                                                                                                                                                                                                                                                                                c                               V       f��     �   /   1  `                  Q <= ;5��    /                     �                     5�_�  �             �   0       ����                                                                                                                                                                                                                                                                                                                c                               V       f��     �   /   1  `                  Q <= D;5��    /                     �                     5�_�  �                0       ����                                                                                                                                                                                                                                                                                                                c                               V       f��     �   /   1  `                  Q <= D();5��    /                  	   �              	       �    /                    �                    5�_�                  0        ����                                                                                                                                                                                                                                                                                                                c                               V       f��     �   /   1  `      !            Q <= D(479 downto 0);5��    /                      �                     5�_�                 0       ����                                                                                                                                                                                                                                                                                                                c                               V       f�f     �   0   2  `    5��    0                      �                     5�_�                 1       ����                                                                                                                                                                                                                                                                                                                d                               V       f�g     �   0   2  a                  5��    0                     �                     5�_�                 1       ����                                                                                                                                                                                                                                                                                                                d                               V       f�i     �   0   2  a                  ()5��    0                  
   �              
       5�_�                 1       ����                                                                                                                                                                                                                                                                                                                d                               V       f�l     �   0   2  a                  (3 downto 0)5��    0                     �                     5�_�                 1       ����                                                                                                                                                                                                                                                                                                                d                               V       f��     �   0   1                       (3 downto 0) & 4bits5��    0                      �      !               5�_�                 /       ����                                                                                                                                                                                                                                                                                                                c           /          /   $       v   $    f��     �   .   0  `      *        elsif clk'event and clk = '1' then5��    .                    �                    �    .                     �                     �    .                     �                     �    .                     �                     �    .                     �                     �    .                    �                    �    .                    �                    �    .                    �                    5�_�    	             /       ����                                                                                                                                                                                                                                                                                                                c           /          /   $       v   $    f��     �   .   0  `              elsif rising_edge then5��    .                     �                     5�_�    
          	   /       ����                                                                                                                                                                                                                                                                                                                c           /          /   $       v   $    f��     �   .   0  `               elsif rising_edge() then5��    .                     �                     5�_�  	            
   /       ����                                                                                                                                                                                                                                                                                                                c           /          /   $       v   $    f��     �   .   0  `      #        elsif rising_edge(clk) then5��    .                     �                     5�_�  
               /       ����                                                                                                                                                                                                                                                                                                                c           /          /   $       v   $    f��     �   .   0  a                  �   .   0  `    5��    .                      r              	       �    .                     r                    �    .                    z                    5�_�                 /   	    ����                                                                                                                                                                                                                                                                                                                d           0          0   $       v   $    f��     �   .   /          
        el5��    .                      r                     5�_�                 /   	    ����                                                                                                                                                                                                                                                                                                                c           /          /   $       v   $    f��     �   /   1  a                  �   /   1  `    5��    /                      �              	       �    /                     �                    �    /                     �                     �    /                     �                     �    /                    �                    �    /                    �                    �    /                 	   �             	       5�_�                 0       ����                                                                                                                                                                                                                                                                                                                d           /          /   $       v   $    f��     �   /   1  a                  if enable = 5��    /                     �                     5�_�                 0       ����                                                                                                                                                                                                                                                                                                                d           /          /   $       v   $    f��     �   /   1  a                  if enable = ''5��    /                     �                     5�_�                 0       ����                                                                                                                                                                                                                                                                                                                d           /          /   $       v   $    f��     �   /   2  a                  if enable = '1'5��    /                     �                     �    /                    �                    �    /                    �                    �    /                    �                    �    /                     �                     �    0                     �                    5�_�                 2       ����                                                                                                                                                                                                                                                                                                                e           /          /   $       v   $    f��     �   1   2          (            Q <= D(479 downto 0) & data;5��    1                      �      )               5�_�                 1        ����                                                                                                                                                                                                                                                                                                                d           1          1          V       f��     �   0   2  `    �   1   2  `    �   0   1                          q5��    0                      �                     �    0                      �              )       5�_�                 1       ����                                                                                                                                                                                                                                                                                                                d           1           1   '       V       f��     �   0   2  a      (            Q <= D(479 downto 0) & data;5��    0                     �                     5�_�                 1       ����                                                                                                                                                                                                                                                                                                                d           1           1   '       V       f��     �   1   4  b                      �   1   3  a    5��    1                      �                     �    1                     �                     �    1                     �                    �    1                    �                     �    2                     �                    �    2                                        5�_�                 3       ����                                                                                                                                                                                                                                                                                                                f           1           1   '       V       f��   k �   3   5  d                      �   3   5  c    5��    3                                           �    3                                          �    3                                         �    3                                          5�_�                 r        ����                                                                                                                                                                                                                                                                                                                g                                            f��     �   r   u  e          �   r   t  d    5��    r                      �	                     �    r                      �	                     �    r                     �	                     �    s                     �	                     �    s                     �	                     �    s                     �	                     �    s                     �	                     5�_�                 t       ����                                                                                                                                                                                                                                                                                                                g                                            f��     �   s   t              5��    s                      �	                     5�_�                 s        ����                                                                                                                                                                                                                                                                                                                g           r           l           V        f��     �   s   {  e    �   s   t  e    5��    s                      �	              �       5�_�                 t       ����                                                                                                                                                                                                                                                                                                                g           r           l           V        f��     �   s   u  l          component reg32 is5��    s                    �	                    �    s                     �	                     �    s                     �	                     �    s                    �	                    �    s                    �	                    �    s                    �	                    5�_�                 v       ����                                                                                                                                                                                                                                                                                                                g           r           l           V        f��     �   u   w  l                  rst, clk: in bit;5��    u                     �	                     �    u                    �	                    �    u                    �	                    �    u                    �	                    5�_�                 v       ����                                                                                                                                                                                                                                                                                                                g           r           l           V        f��     �   v   x  m              �   v   x  l    5��    v                      �	                     �    v                     �	                    5�_�                 w        ����                                                                                                                                                                                                                                                                                                                g           w          w          V       f��     �   v   x  l    �   w   x  l    �   v   w                      data5��    v                      �	                     �    v                      �	              *       5�_�                 w       ����                                                                                                                                                                                                                                                                                                                g           w           w   (       V       f��     �   v   x  m      )        data: in bit_vector(31 downto 0);5��    v                     �	                     5�_�                �       ����                                                                                                                                                                                                                                                                                                                g           w           w   (       V       f�K     �   �   �  m    �   �   �  m    5��    �                      �              .       5�_�    !              �       ����                                                                                                                                                                                                                                                                                                                g           w           w   (       V       f�M     �   �   �  n      -    signal av: bit_vector(31 downto 0) := h0;5��    �                                         �    �                                         �    �                                         �    �                                         5�_�     "          !   �       ����                                                                                                                                                                                                                                                                                                                g           w           w   (       V       f�[     �   �   �  n      0    signal w_vec: bit_vector(31 downto 0) := h0;5��    �                                        5�_�  !  #          "   �   .    ����                                                                                                                                                                                                                                                                                                                g           w           w   (       V       f�_     �   �   �  n      1    signal w_vec: bit_vector(511 downto 0) := h0;5��    �   .                 #                    5�_�  "  $          #   �       ����                                                                                                                                                                                                                                                                                                                g           w           w   (       V       f�f   l �   �   �  n      0    signal k_const, w_vec, kpw_vec: aux_signals;5��    �                     �                     5�_�  #  %          $   �       ����                                                                                                                                                                                                                                                                                                                g           w           w   (       V       f�k     �   �   �  n    5��    �                      "                     �    �                      "                     5�_�  $  &          %   �       ����                                                                                                                                                                                                                                                                                                                g           w           w   (       V       f�n     �   �   �          0    signal current_kpw: bit_vector(31 downto 0);5��    �                            1               5�_�  %  '          &   �        ����                                                                                                                                                                                                                                                                                                                g           w           w   (       V       f�p   m �   �   �  n    �   �   �  n    5��    �                      "              1       5�_�  &  (          '          ����                                                                                                                                                                                                                                                                                                                g                             V       f��     �               #    w_vec(0)  <= msgi(31 downto 0);   $    w_vec(1)  <= msgi(63 downto 32);   $    w_vec(2)  <= msgi(95 downto 64);   %    w_vec(3)  <= msgi(127 downto 96);   &    w_vec(4)  <= msgi(159 downto 128);   &    w_vec(5)  <= msgi(191 downto 160);   &    w_vec(6)  <= msgi(223 downto 192);   &    w_vec(7)  <= msgi(255 downto 224);   &    w_vec(8)  <= msgi(287 downto 256);   &    w_vec(9)  <= msgi(319 downto 288);   &    w_vec(10) <= msgi(351 downto 320);   &    w_vec(11) <= msgi(383 downto 352);   &    w_vec(12) <= msgi(415 downto 384);   &    w_vec(13) <= msgi(447 downto 416);   &    w_vec(14) <= msgi(479 downto 448);   &    w_vec(15) <= msgi(511 downto 480);5��                          o      h              5�_�  '  )          (          ����                                                                                                                                                                                                                                                                                                                g                             V       f��     �                5��                          o                     5�_�  (  *          )  F       ����                                                                                                                                                                                                                                                                                                                g                             V       f�     �  E  G  _                  �  E  G  ^    5��    E                     S$                     �    E                    _$                     5�_�  )  +          *     	    ����                                                                                                                                                                                                                                                                                                                g                             V       f��     �      _      1        	make1: sigma1 port map(w_vec(i-2), op1);5��      	                 �                    5�_�  *  ,          +     	    ����                                                                                                                                                                                                                                                                                                                g                             V       f��     �      _      2        	make2: sigma0 port map(w_vec(i-15), op2);5��      	                                     5�_�  +  -          ,     	    ����                                                                                                                                                                                                                                                                                                                g                             V       f�     �      _      7        	make3: adder32 port map(op3, w_vec(i-7), op3);5��      	                 J                    5�_�  ,  .          -  
       ����                                                                                                                                                                                                                                                                                                                g                             V       f�     �  
    _    5��    
                                          �    
                                          5�_�  -  /          .          ����                                                                                                                                                                                                                                                                                                                g                             V       f�     �      `    �      `    5��                                       �       5�_�  .  0          /     	    ����                                                                                                                                                                                                                                                                                                                g             	         	              f�     �      c      0        	int1: sigma1 port map(w_vec(i-2), op1);5��                                             5�_�  /  1          0     	    ����                                                                                                                                                                                                                                                                                                                g             	         	              f�     �      c      1        	int2: sigma0 port map(w_vec(i-15), op2);5��                        ?                     5�_�  0  2          1     	    ����                                                                                                                                                                                                                                                                                                                g             	         	              f�     �      c      6        	int3: adder32 port map(op3, w_vec(i-7), op3);5��                        l                     5�_�  1  3          2         ����                                                                                                                                                                                                                                                                                                                g             	         	              f�,     �      c    �      c    5��                         �              2       5�_�  2  5          3         ����                                                                                                                                                                                                                                                                                                                g             	         	              f�,     �      d    �      d    5��                         �              2       5�_�  3  6  4      5         ����                                                                                                                                                                                                                                                                                                                g             	         	              f�<     �      e      1    int3: adder32 port map(op3, w_vec(i-7), op3);5��                       �                    5�_�  5  9          6         ����                                                                                                                                                                                                                                                                                                                g             	         	              f�=     �      e      1    int3: adder32 port map(op3, w_vec(i-7), op3);5��                       �                    5�_�  6  :  7      9          ����                                                                                                                                                                                                                                                                                                                g             	         	              f��     �      e      +    int1: sigma1 port map(w_vec(i-2), op1);5��                        /                    5�_�  9  ;          :          ����                                                                                                                                                                                                                                                                                                                g             	         	              f��     �      e      ,    int2: sigma0 port map(w_vec(i-15), op2);5��                        Z                    5�_�  :  <          ;     &    ����                                                                                                                                                                                                                                                                                                                g             	         	              f��     �      e      1    int3: adder32 port map(op3, w_vec(i-7), op3);5��      &                 �                    5�_�  ;  =          <         ����                                                                                                                                                                                                                                                                                                                g             	         	              f��     �      e      /    int3: adder32 port map(op3, w_vec(0), op3);5��                                           �                        �                     �                        �                     �                        �                     �                                           �                                           �                                           5�_�  <  >          =          ����                                                                                                                                                                                                                                                                                                                g             	         	              f��     �      e      1    int3: adder32 port map(w_vec, w_vec(0), op3);5��                         �                     5�_�  =  ?          >     !    ����                                                                                                                                                                                                                                                                                                                g             	         	              f��     �      e      3    int3: adder32 port map(w_vec(), w_vec(0), op3);5��      !                  �                     5�_�  >  @          ?     !    ����                                                                                                                                                                                                                                                                                                                g             	         	              f��     �      e      6    int3: adder32 port map(w_vec(i-7), w_vec(0), op3);5��      !                 �                    5�_�  ?  A          @     !    ����                                                                                                                                                                                                                                                                                                                g             	         	              f��     �              1    int4: adder32 port map(op3, w_vec(i-7), op3);5��                         �      2               5�_�  @  B          A     !    ����                                                                                                                                                                                                                                                                                                                g             	         	              f��     �      d    �      d    5��                         d              2       5�_�  A  C          B          ����                                                                                                                                                                                                                                                                                                                g             	         	              f��     �      e      1    int4: adder32 port map(op3, w_vec(i-7), op3);5��              
          �      
              5�_�  B  D          C         ����                                                                                                                                                                                                                                                                                                                g             	         	              f��     �      e      *    int4: adder32 port map(op3, op2, op3);5��                       �                    5�_�  C  E          D     /    ����                                                                                                                                                                                                                                                                                                                g             	         	              f��     �      e      4    int3: adder32 port map(w_vec(9), w_vec(0), op3);5��      /                 �                    5�_�  D  F          E          ����                                                                                                                                                                                                                                                                                                                g             	         	              f��     �      e      1    int5: adder32 port map(op3, w_vec(i-7), op3);5��              
          �      
              �                        �                    5�_�  E  G          F     %    ����                                                                                                                                                                                                                                                                                                                g             	         	              f��     �      e      *    int5: adder32 port map(op3, op4, op3);5��      %                 �                    �      '                 �                    5�_�  F  H          G          ����                                                                                                                                                                                                                                                                                                                g                      '       v   '    f��     �      e      *    int1: sigma1 port map(w_vec(14), op1);5��                         /                     5�_�  G  I          H         ����                                                                                                                                                                                                                                                                                                                g                      '       v   '    f�     �      e      (    int1: sigma1 port map(w_vec(), op1);�      e    5��                         /                     5�_�  H  J          I          ����                                                                                                                                                                                                                                                                                                                g                               v        f�     �      e      )    int2: sigma0 port map(w_vec(1), op2);�      e    5��                        d                    5�_�  I  K          J     +    ����                                                                                                                                                                                                                                                                                                                g             +         +       v   +    f�     �      e      4    int3: adder32 port map(w_vec(9), w_vec(0), op4);�      e    5��      +                 �                    5�_�  J  L          K     !    ����                                                                                                                                                                                                                                                                                                                g             !         !       v   !    f�3     �      e      A    int3: adder32 port map(w_vec(9), w_vec(511 downto 480), op4);�      e    5��      !                 �                    5�_�  K  M          L     +    ����                                                                                                                                                                                                                                                                                                                g             !         .       v   !    f�;     �              =    	signal op1, op2, op3, op4, op5: bit_vector(31 downto 0);5��                         �      >               5�_�  L  N          M  
        ����                                                                                                                                                                                                                                                                                                                g             !         .       v   !    f�=     �  
    d    �  
    d    5��    
                     �              >       5�_�  M  O          N         ����                                                                                                                                                                                                                                                                                                                g             !         .       v   !    f�>     �  
    e      =    	signal op1, op2, op3, op4, op5: bit_vector(31 downto 0);5��    
                    �                     5�_�  N  P          O         ����                                                                                                                                                                                                                                                                                                                g          	                   V       f�L     �  
            <    signal op1, op2, op3, op4, op5: bit_vector(31 downto 0);5��    
                     �      =               5�_�  O  Q          P   �        ����                                                                                                                                                                                                                                                                                                                g          	                   V       f�S     �   �   �  d    �   �   �  d    5��    �                      T              =       5�_�  P  R          Q   �   "    ����                                                                                                                                                                                                                                                                                                                g           �          �   !       v   !    f�\     �   �   �  e      <    signal op1, op2, op3, op4, op5: bit_vector(31 downto 0);5��    �   "                  v                     �    �   #                  w                     �    �   "                 v                    5�_�  Q  T          R   �   #    ����                                                                                                                                                                                                                                                                                                                g           �          �   !       v   !    f�_     �   �   �  e      >    signal op1, op2, op3, op4, op5, : bit_vector(31 downto 0);�   �   �  e    5��    �   $                  x                     5�_�  R  U  S      T   �   &    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�s     �   �   �  e      U    signal op1, op2, op3, op4, op5, op1, op2, op3, op4, op5: bit_vector(31 downto 0);5��    �   &                 z                    5�_�  T  V          U   �   +    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�v     �   �   �  e      U    signal op1, op2, op3, op4, op5, op6, op2, op3, op4, op5: bit_vector(31 downto 0);5��    �   +                                     5�_�  U  W          V   �   0    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�y     �   �   �  e      U    signal op1, op2, op3, op4, op5, op6, op7, op3, op4, op5: bit_vector(31 downto 0);5��    �   0                 �                    5�_�  V  X          W   �   5    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�|     �   �   �  e      U    signal op1, op2, op3, op4, op5, op6, op7, op8, op4, op5: bit_vector(31 downto 0);5��    �   5                 �                    5�_�  W  Z          X   �   ;    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�}     �   �   �  e      U    signal op1, op2, op3, op4, op5, op6, op7, op8, op9, op5: bit_vector(31 downto 0);5��    �   :                 �                    5�_�  X  [  Y      Z   �   /    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�N     �   �   �  f          �   �   �  e    5��    �                      "                     �    �                     &                     �    �                     7                     �    �                     6                     �    �                    5                    �    �                     7                     �    �                     6                     �    �                 
   5             
       �    �                     >                     �    �                     =                     �    �                     <                     �    �                     ;                     �    �                     :                     �    �                     9                     �    �                     8                     �    �                     7                     �    �                     6                     �    �                 
   5             
       �    �          
          5      
              �    �                 
   5             
       5�_�  Z  \          [   �       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�W     �   �   �  f          signal next_w: bit_vector5��    �                     ?                     5�_�  [  ]          \   �       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�X     �   �   �  f          signal next_w: bit_vector()5��    �                     @                     �    �   %                 G                    5�_�  \  ^          ]   �   *    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�[     �   �   �  f      *    signal next_w: bit_vector(31 downto 0)5��    �   *                  L                     �    �   ,                  N                     �    �   +                  M                     �    �   *                 L                    5�_�  ]  _          ^     %    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�h     �      f      *    int5: adder32 port map(op3, op4, op5);5��      %                 _                    �      '                  a                     �      &                  `                     �      %                 _                    �      %                 _                    �      %                 _                    5�_�  ^  `          _   �   *    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f��     �   �   �  f    �   �   �  f    5��    �                      N              1       5�_�  _  a          `   �       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f��     �   �   �  g      0    signal current_kpw: bit_vector(31 downto 0);5��    �                    a                    5�_�  `  b          a         ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f��     �      h          �      g    5��                         �                     �                        �                     �                        �                     �                        �                     �                        �                     �                        �                     �                    	   �             	       �             	          �      	              �                    	   �             	       5�_�  a  c          b         ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f��     �      h          current_w5��                        �                     �                        �                     �                       �                    �                       �                    �                       �                    5�_�  b  d          c         ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f��     �      h          current_w <= w_vec5��                        �                     5�_�  c  e          d         ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f��     �      h          current_w <= w_vec()5��                        �                     5�_�  d  f          e     &    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f��     �      h      &    current_w <= w_vec(511 downto 480)5��      &                  �                     5�_�  e  g          f     &    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�     �      i          �      h    5��                         �                     �                        �                     5�_�  f  h          g         ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�(     �      j          �      i    5��                         �                     �                        �                     �                    	   �             	       �                        �                     �                       �                    �                        �                     �                        �                     �                        �                     �                        �                     �                       �                    �                       �                    �                       �                    �                        �                     �                       �                    �                       �                    �                    	   �             	       5�_�  g  i          h     !    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�;     �      j      !    shf_w: shift_reg512 port map 5��      !                  �                     5�_�  h  j          i     "    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�?     �      j      #    shf_w: shift_reg512 port map ()5��      "                  �                     5�_�  i  k          j     "    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�S     �      j      &    shf_w: shift_reg512 port map (clk)5��      "                  �                     5�_�  j  l          k     *    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�V     �      j      +    shf_w: shift_reg512 port map (rst, clk)5��      *                  �                     �      ,                  �                     �      +                 �                    5�_�  k  m          l     ,    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�Z     �      j      -    shf_w: shift_reg512 port map (rst, clk, )5��      ,                  �                     5�_�  l  n          m     -    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�[     �      j      /    shf_w: shift_reg512 port map (rst, clk, '')5��      -                                        5�_�  m  o          n     /    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�]   n �      j      0    shf_w: shift_reg512 port map (rst, clk, '1')5��      /                                       5�_�  n  p          o   �   -    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�     �   �   �  j    �   �   �  j    5��    �                      }              /       5�_�  o  q          p   �       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�     �   �   �  k      .    signal current_w: bit_vector(31 downto 0);5��    �                    �                    5�_�  p  r          q         ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�1     �     "  m          get_kpw: adder32�    "  l              �    !  k    5��                         =               	       �                         =                      �                        =               	       �                        B                     �                        K                     �                        K                     �                        K                     5�_�  q  s          r  !       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�\     �     "  m          get_kpw: adder325��                         R                      �                        S                     �                        S                     �                     	   S              	       5�_�  r  t          s  !       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�a     �     "  m          get_kpw: adder32 port map 5��                         \                      5�_�  s  u          t  !       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�e     �     "  m           get_kpw: adder32 port map ()5��                         ]                      �                     	   ]              	       �              	          ]       	              �                        ]                     �       *              	   h              	       �       *       	          h       	              �       *              	   h              	       �       2                 p                     5�_�  t  v          u  !   3    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�k     �     "  m      4    get_kpw: adder32 port map (current_w, current_k)5��       3                  q                      �       5                 s                     �       5                 s                     �       5                 s                     �       5                 s                     5�_�  u  w          v  !   A    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�o     �     "  m      A    get_kpw: adder32 port map (current_w, current_k, current_kpw)5��       A                                        5�_�  v  x          w  T       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�     �  S  U  m                  -- Calculate W5��    S                
   �&             
       5�_�  w  y          x  U       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�&     �  T  V  n                  �  T  V  m    5��    T                     �&                     �    T                    �&                     �    T                   �&                    �    T                	   �&             	       �    T         	       	   �&      	       	       �    T         	          �&      	              �    T                
   �&             
       �    T                   �&                    �    T                   �&                    �    T                   �&                    �    T                   �&                    �    T                   �&                    5�_�  x  z          y  U        ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�;     �  T  V  n                   current_k <= k_const5��    T                     �&                     5�_�  y  {          z  U   !    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�A     �  T  V  n      "            current_k <= k_const()5��    T  !                  �&                     �    T  !              	   �&             	       �    T  !       	          �&      	              �    T  !              	   �&             	       5�_�  z  |          {  U   +    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�D     �  T  V  n      +            current_k <= k_const(iteration)5��    T  +                   '                     5�_�  {  }          |  U   +    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�<     �  U  W  n    �  U  V  n    5��    U                     '              -       5�_�  |  ~          }  V       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�@     �  U  W  o      ,            current_k <= k_const(iteration);5��    U                   '                    5�_�  }            ~  V       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�G     �  U  W  o      ,            current_w <= k_const(iteration);5��    U                   '                    5�_�  ~  �            V       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�K     �  U  W  o      &            current_w <= w(iteration);5��    U                    '                     �    U                   '                    �    U                   '                    �    U                   '                    5�_�    �          �  V       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�M   o �  U  W  o      *            current_w <= w_vec(iteration);5��    U         	          !'      	              �    U  #                 %'                    �    U  #                 %'                    �    U  #              
   %'             
       5�_�  �  �          �  W   ,    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�]     �  V  W          .            current_kpw <= kpw_vec(iteration);5��    V                     2'      /               5�_�  �  �  �      �         ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f��     �              '    current_w <= w_vec(511 downto 480);5��                         �      (               5�_�  �  �          �     1    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f��     �      m      2    shf_w: shift_reg512 port map (rst, clk, '1', )5��      1                                       �      1                                     �      1                                     �      1                                     5�_�  �  �          �     7    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f��     �      m      8    shf_w: shift_reg512 port map (rst, clk, '1', next_w)5��      7                                       5�_�  �  �          �     +    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�     �      m      :    shf_w: shift_reg512 port map (rst, clk, '1', next_w, )5��      +                                       5�_�  �  �          �     +    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�     �      m      6    shf_w: shift_reg512 port map (rst, clk,, next_w, )5��      +                                       5�_�  �  �          �     4    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�     �      m      5    shf_w: shift_reg512 port map (rst, clk, next_w, )5��      4                                       �      4                                     �      4                                     �      4                                     5�_�  �  �          �     :    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�7     �      m      :    shf_w: shift_reg512 port map (rst, clk, next_w, w_vec)5��      :                                       5�_�  �  �          �   v       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�?     �   u   w  m      %            rst, clk, enable: in bit;5��    u                     �	                     5�_�  �  �          �   (       ����                                                                                                                                                                                                                                                                                                                g           E   (       E          v       f��     �   '   )  m          �   (   )  m    5��    '                  %   	              %       5�_�  �  �          �   (   '    ����                                                                                                                                                                                                                                                                                                                g           E   (       E          v       f��     �   (   *  m    5��    (                      0                     �    (                      0                     5�_�  �  �          �   (   
    ����                                                                                                                                                                                                                                                                                                                h           F   (       F          v       f��     �   '   )  n      )   signal counter: unsigned(5 downto 0); 5��    '   
                                     5�_�  �  �          �   (       ����                                                                                                                                                                                                                                                                                                                h           F   (       F          v       f��     �   '   )  n      (   signal vector: unsigned(5 downto 0); 5��    '                                        �    '                                          �    '                                          �    '                                          �    '                 
                
       �    '          
                
              �    '                 
                
       5�_�  �  �          �   (       ����                                                                                                                                                                                                                                                                                                                h           F   (       F          v       f��     �   '   )  n      *   signal vector: bit_vector(5 downto 0); 5��    '                     $                     5�_�  �  �  �      �   1       ����                                                                                                                                                                                                                                                                                                                h           F   (       F          v       f�     �   0   1                       if enable = '1' then5��    0                      �      !               5�_�  �  �          �   2       ����                                                                                                                                                                                                                                                                                                                g           E   (       E          v       f�     �   1   2                      else                   Q <= D;5��    1                      �      )               5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                e           C   (       C          v       f�      �   0   2  k      ,                Q <= D(479 downto 0) & data;5��    0                     �                     5�_�  �  �          �   2       ����                                                                                                                                                                                                                                                                                                                e           C   (       C          v       f�!     �   1   2                      end if;5��    1                      �                     5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                d           B   (       B          v       f�,     �   0   2  j      (            Q <= D(479 downto 0) & data;5��    0                    �                    �    0                     �                     �    0                     �                     �    0                    �                    �    0                    �                    �    0                    �                    5�_�  �  �          �   3       ����                                                                                                                                                                                                                                                                                                                d           B   (       B          v       f�D     �   4   6  l          Q <= vector�   3   6  k          �   3   5  j    5��    3                                           �    3                                           �    3                                          �    4                                          �    4                                          �    4   
                                       �    4   	                                     �    4   	                                     �    4   	                                     5�_�  �  �          �   /       ����                                                                                                                                                                                                                                                                                                                f           /          /          v       f��     �   .   0  l      !            Q <= (others => '0');5��    .                    �                    5�_�  �  �          �   /       ����                                                                                                                                                                                                                                                                                                                f           /          /          v       f��     �   .   0  l                  Q <= d;5��    .                    �                    5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                f           /          /          v       f��     �   0   2  l      -            Q <= vector(479 downto 0) & data;5��    0                    �                    5�_�  �  �          �   5       ����                                                                                                                                                                                                                                                                                                                f           /          /          v       f��     �   4   6  l          Q <= vector;5��    4                                        5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                f           /          /          v       f��     �      !  l      !        rst, clk, enable: in bit;5��                         0                     5�_�  �  �          �     3    ����                                                                                                                                                                                                                                                                                                                f           /          /          v       f �     �      l      ;    shf_w: shift_reg512 port map (rst, clk, next_w, w_vec);5��      3                  �                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                f           /          /          v       f �     �           
   %    get_w: for i in 16 to 63 generate   
    	begin   0        	int1: sigma1 port map(w_vec(i-2), op1);   1        	int2: sigma0 port map(w_vec(i-15), op2);   6        	int3: adder32 port map(op3, w_vec(i-7), op3);   0        	make4: adder32 port map(op3, op2, op4);   8        	make5: adder32 port map(op4, w_vec(i-16), op5);           	w_vec(i) <= op5;       end generate;    5��          
                     b              5�_�  �  �          �     4    ����                                                                                                                                                                                                                                                                                                                f           /          /          v       f �     �      b      4    int1: sigma1 port map(w_vec(63 downto 32), op1);5��      4                  X                     5�_�  �  �          �     8    ����                                                                                                                                                                                                                                                                                                                f           /          /          v       f �     �      b      8    int1: sigma1 port map(w_vec(63 downto 32), op1); -- 5��      8                  \                     5�_�  �  �          �     6    ����                                                                                                                                                                                                                                                                                                                f           /          /          v       f �     �      b      6    int2: sigma0 port map(w_vec(479 downto 448), op2);5��      6                  �                     5�_�  �  �          �     N    ����                                                                                                                                                                                                                                                                                                                f           /          /          v       f �     �    	  b      N    int3: adder32 port map(w_vec(223 downto 192), w_vec(511 downto 480), op4);5��      N                                       5�_�  �  �          �     R    ����                                                                                                                                                                                                                                                                                                                f           /          /          v       f �     �    	  b      R    int3: adder32 port map(w_vec(223 downto 192), w_vec(511 downto 480), op4); -- 5��      R               
                 
       5�_�  �  �          �     \    ����                                                                                                                                                                                                                                                                                                                f           /          /          v       f �     �    	  b      \    int3: adder32 port map(w_vec(223 downto 192), w_vec(511 downto 480), op4); -- t-9 and t-5��      [                  %                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    f �     �              (    get_kpw: for j in 0 to 63 generate     3    	signal op1, op2, op3: bit_vector(31 downto 0);           begin           	op1 <= w_vec(j);               op2 <= k_const(j);   0        	make1: adder32 port map(op1, op2, op3);               kpw_vec(j) <= op3;       	end generate;5��                         �                    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    f �   q �               5��                         �                     5�_�  �  �          �   w       ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fqe     �   v   x  Y      *            d: in bit_vector(31 downto 0);5��    v                    �	                    5�_�  �  �          �   x       ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fqi   r �   w   y  Y      *            q: out bit_vector(31 downto 0)5��    w                    
                    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    frZ     �   �   �  Y      )    signal k_const, kpw_vec: aux_signals;5��    �                     u                     5�_�  �  �  �      �   �       ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fr]     �   �   �  Y      "    signal k_const, : aux_signals;5��    �                     s                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    frf     �   �   �  Y      V    signal op1, op2, op3, op4, op5, op6, op7, op8, op9, op10: bit_vector(31 downto 0);5��    �                     �                     5�_�  �  �          �  A   +    ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fr�   s �  @  B  Y      /            current_w <= w_vec(511 downto 479);5��    @  +                 `$                    5�_�  �  �          �  
   8    ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fr�     �      [          get_w: reg32 port�  
    Z          �  
    Y    5��    
                     p                     �    
                    t                     �    
                    t                     �    
                   t                     �                        y                     �                       |                    �                        �                     �                        �                     �                       �                    �                       �                    �                    	   �             	       5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fs     �      [          get_w: reg32 port map 5��                        �                     5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fs     �      [          get_w: reg32 port map ()5��                     	   �              	       �      #                 �                    �      %                 �                    �      %                 �                    �      %                 �                    5�_�  �  �          �     *    ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fs     �      [      +    get_w: reg32 port map (rst, clk, w_vec)5��      *                  �                     5�_�  �  �          �     +    ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fs     �      [      -    get_w: reg32 port map (rst, clk, w_vec())5��      +                  �                     �      /                 �                    �      /                 �                    �      /              
   �             
       5�_�  �  �          �     :    ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fs     �      [      ;    get_w: reg32 port map (rst, clk, w_vec(511 downto 480))5��      :                  �                     �      <              	   �             	       �      <       	          �      	              �      <              	   �             	       5�_�  �  �          �     F    ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fs      �      [      F    get_w: reg32 port map (rst, clk, w_vec(511 downto 480), current_w)5��      F                  �                     5�_�  �  �  �      �  C   .    ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    ft�     �  B  C          /            current_w <= w_vec(511 downto 480);5��    B                     �$      0               5�_�  �  �          �   �   *    ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    ft�   w �   �   �  Z      3    signal w_vec: bit_vector(511 downto 0) := msgi;5��    �   *                  �                     5�_�  �  �          �  B   %    ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fv�     �  B  D  [                  �  B  D  Z    5��    B                     z$                     �    B                    �$                     �    B                    �$                     �    B                    �$                     �    B                	   �$             	       �    B         	          �$      	              �    B                   �$                    5�_�  �  �          �  C       ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fv�     �  B  D  [                  current_w <= �  C  D  [    5��    B                    �$                     5�_�  �  �          �  C   .    ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fv�     �  B  D  [      .            current_w <= w_vec(511 downto 480)5��    B  .                  �$                     5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fv�     �  
                   G    get_w: reg32 port map (rst, clk, w_vec(511 downto 480), current_w);5��    
                     h      M               5�_�  �  �  �      �  
        ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fv�     �  	    Y    5��    	                     &                     �    	                     &                     5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fw     �      Z          -- W iterations5��                        �                     �      	                 �                    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fw     �  
    [          �  
    Z    5��    
                     *                     �    
                    .                     5�_�  �  �          �   (   *    ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fw�     �   '   )  [      ,   signal vector: bit_vector(511 downto 0); 5��    '   *                  (                     5�_�  �  �          �   /       ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fw�     �   .   0  [                  q <= d;5��    .                    �                    �    .                     �                     �    .                     �                     �    .                     �                     �    .                    �                    �    .                    �                    �    .                    �                    5�_�  �  �          �   /       ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fw�     �   .   0  [                  vector <= d5��    .                     �                     5�_�  �  �          �   (   *    ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fw�   x �   '   )  [      1   signal vector: bit_vector(511 downto 0) := d; 5��    '   *                  (                     5�_�  �  �          �   �   *    ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fw�     �   �   �  [      +    signal w_vec: bit_vector(511 downto 0);5��    �   *                  �                     �    �   0                 �                    5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fx      �   0   2  [      -            q <= vector(479 downto 0) & data;5��    0                    �                    5�_�  �  �          �   �   *    ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fx.   y �   �   �  [      3    signal w_vec: bit_vector(511 downto 0) := msgi;5��    �   *                  �                     5�_�  �  �          �  ;       ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fz   z �  ;  =  \                  �  ;  =  [    5��    ;                     �#                     �    ;                    �#                     �    ;                   �#                    �    ;                   �#                    �    ;                   �#                    �    ;                    �#                     �    ;                   �#                    �    ;                   �#                    �    ;                   �#                    5�_�  �  �          �   .       ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fzY   { �   -   /  \              if rst = '0' then5��    -                    i                    5�_�  �  �          �  <       ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fz|   | �  ;  <                      w_vec <= msgi;5��    ;                     �#                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                f                        $       v   $    f}G     �        [      *        elsif clk'event and clk = '1' then5��                        b                    �                         d                     �                        c                    �                         f                     �                         e                     �                         d                     �                         c                     �                        b                    �                        b                    �                        b                    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                f                        $       v   $    f}K     �        [              elsif rising_edge then5��                         m                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                f                        $       v   $    f}K   } �        [               elsif rising_edge() then5��                         n                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                f                        $       v   $    f}�     �        \          �        [    5��                          ^               	       �                         ^                     �                     
   o              
       �              
          o       
              �                     
   o              
       5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                g                        $       v   $    f}�     �        \              init: in bit_vector5��                         y                      5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                g                        $       v   $    f}�     �        \              init: in bit_vector()5��                         z                      �                        }                     �                        }                     �                        }                     5�_�  �  �          �      (    ����                                                                                                                                                                                                                                                                                                                g                        $       v   $    f}�     �        \      (        init: in bit_vector(31 downto 0)5��       (                  �                      5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                g                        $       v   $    f}�     �        \          5��                                              �                                              �                                            �                                            �                                            �                                            5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                g                               v       f}�     �        \          signed(7 downto 0)5��                                            �                                              �                                              �                                              �                                            �                                            �                                            �                         (                     �                         '                     �                        &                    �                         (                     �                         '                     �                     
   &             
       �                         /                     �                         .                     �                         -                     �                         ,                     �                         +                     �                         *                     �                         )                     �                         (                     �                         '                     �                     
   &             
       �              
          &      
              �                     
   &             
       5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                g                               v       f}�     �        \          signal initial: bit_vector5��                         0                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                g                               v       f}�     �        \           signal initial: bit_vector()5��                         1                     �                          2                     �                        1                    �       %                  7                     �       $                  6                     �       #                  5                     �       "                 4                    �       "                 4                    �       "                 4                    5�_�  �  �          �      +    ����                                                                                                                                                                                                                                                                                                                g                               v       f}�     �        \      +    signal initial: bit_vector(31 downto 0)5��       +                  =                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                g                               v       f}�     �        \      !            Q <= (others => '0');5��                         �                     �                         �                     �                        �                    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                g                               v       f}�     �        \                  Q <= init;5��                        �                    �                         �                     �                         �                     �                        �                    �                         �                     �                         �                     �                         �                     �                        �                    �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                g                               v       f}�     �        \                  Q <= D;5��                        �                    �                         �                     �                         �                     �                         �                     �                        �                    �                         �                     �                         �                     �                         �                     �                        �                    �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                g                               v       f}�     �        ]          �        \    5��                                                �                                                �                                               �                                              5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                i                               v       f}�     �        ^      ,    signal initial: bit_vector(31 downto 0);5��                                            5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                i                               v       f}�     �        ^                  initial <= init;5��                        �                    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                i                               v       f}�     �        ^                  initial <= D;5��                        �                    5�_�  �  �          �      	    ����                                                                                                                                                                                                                                                                                                                i                               v       f}�   ~ �        ^      	    q <= 5��       	                                       5�_�  �  �          �   �   &    ����                                                                                                                                                                                                                                                                                                                i           �   &       �   +          +    f~      �   �   �  ^      -    signal av: bit_vector(31 downto 0) := h0;   -    signal bv: bit_vector(31 downto 0) := h1;   -    signal cv: bit_vector(31 downto 0) := h2;   -    signal dv: bit_vector(31 downto 0) := h3;   -    signal ev: bit_vector(31 downto 0) := h4;   -    signal fv: bit_vector(31 downto 0) := h5;   -    signal gv: bit_vector(31 downto 0) := h6;   -    signal hv: bit_vector(31 downto 0) := h7;5��    �   &                  N                     �    �   &                  v                     �    �   &                  �                     �    �   &                  �                     �    �   &                  �                     �    �   &                                       �    �   &                  >                     �    �   &                  f                     5�_�  �  �          �   �   )    ����                                                                                                                                                                                                                                                                                                                i           �   )       �   .          .    f~(     �   �   �  ^      0    signal a_reg: bit_vector(31 downto 0) := h0;   0    signal b_reg: bit_vector(31 downto 0) := h1;   0    signal c_reg: bit_vector(31 downto 0) := h2;   0    signal d_reg: bit_vector(31 downto 0) := h3;   0    signal e_reg: bit_vector(31 downto 0) := h4;   0    signal f_reg: bit_vector(31 downto 0) := h5;   0    signal g_reg: bit_vector(31 downto 0) := h6;   0    signal h_reg: bit_vector(31 downto 0) := h7;5��    �   )                  �                     �    �   )                  �                     �    �   )                  �                     �    �   )                                       �    �   )                  =                     �    �   )                  h                     �    �   )                  �                     �    �   )                  �                     5�_�  �  �          �     )    ����                                                                                                                                                                                                                                                                                                                i             )         )          )    f~7     �      ^      5    b_register: reg32 port map (rst, clk, bv, b_reg);   5    c_register: reg32 port map (rst, clk, cv, c_reg);   5    d_register: reg32 port map (rst, clk, dv, d_reg);   5    e_register: reg32 port map (rst, clk, ev, e_reg);   5    f_register: reg32 port map (rst, clk, fv, f_reg);   5    g_register: reg32 port map (rst, clk, gv, g_reg);   5    h_register: reg32 port map (rst, clk, hv, h_reg);�      ^      5    a_register: reg32 port map (rst, clk, av, a_reg);5��      )                  *                     �      )                  d                     �      )                  �                     �      )                  �                     �      )                                       �      )                  L                     �      )                  �                     �      )                  �                     5�_�  �  �          �     +    ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f~I     �      ^      9    b_register: reg32 port map (rst, clk, h0, bv, b_reg);   9    c_register: reg32 port map (rst, clk, h0, cv, c_reg);   9    d_register: reg32 port map (rst, clk, h0, dv, d_reg);   9    e_register: reg32 port map (rst, clk, h0, ev, e_reg);   9    f_register: reg32 port map (rst, clk, h0, fv, f_reg);   9    g_register: reg32 port map (rst, clk, h0, gv, g_reg);   9    h_register: reg32 port map (rst, clk, h0, hv, h_reg);5��      +                 f                    �      +                 �                    �      +                 �                    �      +                                     �      +                 N                    �      +                 �                    �      +                 �                    5�_�  �  �  �      �   p       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f~U     �   p   r  _              �   p   r  ^    5��    p                      E	                     �    p                     E	                    �    p                     R	                     �    p                    Q	                    �    p                     \	                     �    p                     [	                     �    p                    Z	                    �    p                     \	                     �    p                     [	                     �    p                 
   Z	             
       �    p                     c	                     �    p                     b	                     �    p                     a	                     �    p                     `	                     �    p                     _	                     �    p                     ^	                     �    p                     ]	                     �    p                     \	                     �    p                     [	                     �    p                 
   Z	             
       �    p          
          Z	      
              �    p                 
   Z	             
       5�_�  �  �          �   q       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f~`     �   p   r  _                  init: in bit_vector5��    p                     d	                     5�_�  �  �          �   q        ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f~`     �   p   r  _      !            init: in bit_vector()5��    p                      e	                     �    p   %                  j	                     �    p   $                  i	                     �    p   #                 h	                    �    p   #                 h	                    �    p   #                 h	                    5�_�  �  �          �   q   ,    ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f~c    �   p   r  _      ,            init: in bit_vector(31 downto 0)5��    p   ,                  q	                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f$   � �        _              if rst = '0' then5��                        z                    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�     �        _              rst, clk: in bit;5��                         T                      5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�     �        `              �        _    5��                          p                     �                         p                    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                j             +         +          +    f�     �                        if ena5��                          p                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�     �        `              �        _    5��                          p              	       �                         x                     �                         }                     �                         |                     �                        {                    �                        {                    �                        {                    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                j             +         +          +    f�     �                        if enable5��                          p                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�     �        _      #        elsif rising_edge(clk) then5��                         �                     �       %                  �                     �       $                  �                     �       #                 �                    �       #                 �                    �       #              	   �             	       �       +                 �                    �       ,                  �                     5�_�  �  �          �      ,    ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�     �        _      1        elsif rising_edge(clk) and enable =  then5��       ,                  �                     5�_�  �  �          �      -    ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�     �        _      3        elsif rising_edge(clk) and enable = '' then5��       -                  �                     5�_�  �  �          �   #       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�3     �   "   $  _              rst, clk: in bit;5��    "                     �                     5�_�  �  �          �   3       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�>     �   2   4  _      $        elsif rising_edge(clk)  then5��    2                     !                     �    2   %                  '                     �    2   $                  &                     �    2   #                 %                    �    2   #                 %                    �    2   #              	   %             	       5�_�  �  �          �   3   ,    ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�A     �   2   4  _      1        elsif rising_edge(clk) and enable =  then5��    2   ,                  .                     5�_�  �  �          �   3   -    ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�C     �   2   4  _      3        elsif rising_edge(clk) and enable = '' then5��    2   -                  /                     5�_�  �  �          �   A       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�R     �   @   B  _      C        clk, rst: in bit;                            -- Clock input5��    @                                          �    @                                          �    @                                          �    @                                        �    @                                        �    @                                        5�_�  �  �          �   O       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�Y     �   N   P  _      #        elsif rising_edge(clk) then5��    N                     �                     �    N   #                 �                    5�_�  �  �          �   �   "    ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�x     �   �   �  `          �   �   �  _    5��    �                      �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    �    �                     �                     �    �                     �                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f��     �   �   �  `          signal enable: bit := 5��    �                     �                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f��     �   �   �  `          signal enable: bit := ""5��    �                     �                     �    �                    �                    �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    5�_�  �  �          �  @       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f��     �  @  B  a                  �  @  B  `    5��    @                     A$                     �    @                    M$                     �    @                    O$                     �    @                    N$                     �    @                   M$                    �    @                   M$                    �    @                
   M$             
       5�_�  �             �  A       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f��     �  @  B  a                  enable <= 5��    @                    W$                     5�_�  �               A       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f��     �  @  B  a                  enable <= ''5��    @                    X$                     5�_�                 A       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f��     �  @  B  a                  enable <= '1'5��    @                    Z$                     5�_�                A       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f��     �  @  B  a                  enable <= '1';5��    @                   X$                    5�_�                ?       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�     �  >  @  b              �  >  @  a    5��    >                     $              	       �    >                    $                     �    >                    $                     �    >                   $                    �    >                   $                    �    >                   $                    5�_�                ?       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�     �  >  @  b              if rst = 5��    >                    $                     5�_�                ?       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�     �  >  @  b              if rst = ''5��    >                     $                     5�_�                ?       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�     �  ?  A  c                  enable�  >  A  b              if rst = '0'5��    >                    "$                     �    >                    '$                     �    >                   '$              	       �    ?                    ($                    �    ?                    6$                     �    ?                    5$                     �    ?                   4$                    �    ?                   4$                    �    ?                	   4$             	       5�_�                @       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�     �  ?  A  c                  enable = 5��    ?                    =$                     5�_�    	            @       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�     �  ?  A  c                  enable = ''5��    ?                    >$                     �    ?                   >$                    5�_�    
          	  @       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�     �  ?  B  c                  enable = '1'5��    ?                    @$                     �    ?                   A$                     �    @                    N$                     �    @                    B$                    �    @                    N$                     5�_�  	            
  @       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�   � �  ?  A  d                  enable = '1';5��    ?                    ;$                     5�_�  
               *    ����                                                                                                                                                                                                                                                                                                                i             )         )          )    f�;     �      d      9    b_register: reg32 port map (rst, clk, h1, bv, b_reg);   9    c_register: reg32 port map (rst, clk, h2, cv, c_reg);   9    d_register: reg32 port map (rst, clk, h3, dv, d_reg);   9    e_register: reg32 port map (rst, clk, h4, ev, e_reg);   9    f_register: reg32 port map (rst, clk, h5, fv, f_reg);   9    g_register: reg32 port map (rst, clk, h6, gv, g_reg);   9    h_register: reg32 port map (rst, clk, h7, hv, h_reg);�      d      9    a_register: reg32 port map (rst, clk, h0, av, a_reg);5��      *                  �                     �      *                                       �      *                  J                     �      *                  �                     �      *                  �                     �      *                                        �      *                  R                      �      *                  �                      5�_�                   -    ����                                                                                                                                                                                                                                                                                                                i             )         )          )    f�C     �      d      9    counter: counter_6bit port map (clk, rst, iteration);5��      -                  �                     �      0                  �                     �      /                  �                     �      .                 �                    �      .                 �                    �      .                 �                    5�_�                   +    ����                                                                                                                                                                                                                                                                                                                i             )         )          )    f�J     �      d      A    shf_w: shift_reg512 port map (rst, clk, next_w, msgi, w_vec);5��      +                                       �      .                                       �      -                                       �      ,                                     �      ,                                     �      ,                                     5�_�                 �       ����                                                                                                                                                                                                                                                                                                                i             )         )          )    f�X     �   �   �  d      G            clk, rst: in bit;                            -- Clock input5��    �                     d                     5�_�                 y       ����                                                                                                                                                                                                                                                                                                                i             )         )          )    f�\     �   x   z  d                  rst, clk: in bit;5��    x                     s
                     5�_�                 p       ����                                                                                                                                                                                                                                                                                                                i             )         )          )    f�d   � �   o   q  d                  rst, clk: in bit;5��    o                     �	                     5�_�                       ����                                                                                                                                                                                                                                                                                                                i             )         )          )    f�     �      f          get_k: reg32�      e          �      d    5��                         �                     �                         �                     �                        �                     �                     
   �              
       �                        �                     �                        �                     �                       �                    �                       �                    �                       �                    �                        �                     �                       �                    �                       �                    �                    	   �             	       5�_�                       ����                                                                                                                                                                                                                                                                                                                i              )         )          )    f�#     �      f          get_k: reg32 port map 5��                        �                     5�_�                       ����                                                                                                                                                                                                                                                                                                                i              )         )          )    f�&     �      f          get_k: reg32 port map ()5��                     	   �              	       �      #                 �                    �      '                  �                     �      &                  �                     �      %                 �                    �      %                 �                    �      %              
   �             
       �      .                  �                     5�_�                   .    ����                                                                                                                                                                                                                                                                                                                i              )         )          )    f�7     �      f      /    get_k: reg32 port map (rst, clk, enable, k)5��      .                  �                     5�_�                   /    ����                                                                                                                                                                                                                                                                                                                i              )         )          )    f�7     �      f      1    get_k: reg32 port map (rst, clk, enable, k())5��      /                  �                     5�_�                   1    ����                                                                                                                                                                                                                                                                                                                i              )         )          )    f�9     �      f      2    get_k: reg32 port map (rst, clk, enable, k(0))5��      1                  �                     �      =                                       �      <                                        �      ;              	   �             	       �      ;       	          �      	              �      ;              	   �             	       �      C                                     5�_�                   E    ����                                                                                                                                                                                                                                                                                                                i              )         )          )    f�x     �      f      E    get_k: reg32 port map (rst, clk, enable, k(0), next_k, current_k)5��      E                  	                     5�_�                   .    ����                                                                                                                                                                                                                                                                                                                i              )         )          )    f��     �      f      F    get_k: reg32 port map (rst, clk, enable, k(0), next_k, current_k);5��      .                  �                     5�_�                 �   *    ����                                                                                                                                                                                                                                                                                                                i              )         )          )    f��     �   �   �  f    �   �   �  f    5��    �                                    ,       5�_�                 �       ����                                                                                                                                                                                                                                                                                                                i          !   )         )          )    f��     �   �   �  g      +    signal next_w: bit_vector(31 downto 0);5��    �                    #                    5�_�                N   *    ����                                                                                                                                                                                                                                                                                                                i          !   )         )          )    f��   � �  M  O  g      ,            current_k <= k_const(iteration);5��    M  *                  @&                     �    M  *                 @&                    5�_�                N       ����                                                                                                                                                                                                                                                                                                                i          !   )         )          )    f��   � �  M  O  g      .            current_k <= k_const(iteration+1);5��    M         	          "&      	              �    M                    #&                     �    M                   "&                    �    M                    '&                     �    M                    &&                     �    M                    %&                     �    M                    $&                     �    M                    #&                     �    M                   "&                    �    M                    '&                     �    M                    &&                     �    M                    %&                     �    M                    $&                     �    M                    #&                     �    M                   "&                    �    M                   "&                    �    M                   "&                    5�_�                M       ����                                                                                                                                                                                                                                                                                                                i          !   )         )          )    f��     �  M  O  h                  �  M  O  g    5��    M                     &                     �    M                    "&                     �    M                   #&                    �    M                    '&                     �    M                    &&                     �    M                	   %&             	       �    M         	          %&      	              �    M                   %&                    5�_�                 O       ����                                                                                                                                                                                                                                                                                                                i          !   )         )          )    f��     �  N  P  h      +            next_k <= k_const(iteration+1);5��    N                    E&                     5�_�    !             O       ����                                                                                                                                                                                                                                                                                                                i          !   )         )          )    f��     �  O  Q  i                      �  O  Q  h    5��    O                     i&                     �    O                    y&                     �    O                    i&                    �    O                    y&                     5�_�     "          !  P       ����                                                                                                                                                                                                                                                                                                                i          !   )         )          )    f��   � �  O  Q  i                  end if.5��    O                   {&                    5�_�  !  #          "  N       ����                                                                                                                                                                                                                                                                                                                i                                            f�     �  M  O  i      "            if iteration < 64 then5��    M                   2&                    5�_�  "  $          #  N       ����                                                                                                                                                                                                                                                                                                                i                                            f�   � �  M  O  i      "            if iteration < 63 then5��    M                   2&                    5�_�  #  &          $  Q       ����                                                                                                                                                                                                                                                                                                                i                                            f��     �  P  Q          /            current_w <= w_vec(511 downto 480);5��    P                     }&      0               5�_�  $  '  %      &  Q       ����                                                                                                                                                                                                                                                                                                                i                                            f��     �  Q  S  h    �  Q  R  h    5��    Q                     �&              0       5�_�  &  (          '  R       ����                                                                                                                                                                                                                                                                                                                i                                            f��     �  Q  S  i      /            current_w <= w_vec(511 downto 480);5��    Q                    �&                     5�_�  '  )          (  R       ����                                                                                                                                                                                                                                                                                                                i                                            f��     �  Q  S  j              �  Q  S  i    5��    Q                     �&              	       �    Q                    �&                     �    Q  
                  �&                     �    Q  	                  �&                     �    Q                	   �&             	       �    Q                    �&                     �    Q                    �&                     �    Q                    �&                     �    Q                    �&                     �    Q                    �&                     �    Q                    �&                     �    Q  
                  �&                     �    Q  	                  �&                     �    Q                	   �&             	       �    Q                    �&                     �    Q                    �&                     �    Q                    �&                     �    Q                    �&                     �    Q                    �&                     �    Q                    �&                     �    Q  
                  �&                     �    Q  	                  �&                     �    Q                	   �&             	       �    Q         	          �&      	              �    Q                   �&                    �    Q                    �&                     �    Q                    �&                     �    Q                   �&                    �    Q                   �&                    �    Q                   �&                    5�_�  (  *          )  R       ����                                                                                                                                                                                                                                                                                                                i                                            f��     �  Q  S  j              current_k <= k_const5��    Q                    �&                     5�_�  )  +          *  R       ����                                                                                                                                                                                                                                                                                                                i                                            f��     �  Q  S  j              current_k <= k_const()5��    Q                    �&                     �    Q                	   �&             	       �    Q         	          �&      	              �    Q                	   �&             	       5�_�  *  ,          +  R   '    ����                                                                                                                                                                                                                                                                                                                i                                            f��     �  Q  S  j      '        current_k <= k_const(iteration)5��    Q  '                  �&                     5�_�  +  -          ,  N   "    ����                                                                                                                                                                                                                                                                                                                i          P         N   "       V   '    f�      �  M  N          "            if iteration < 62 then   /                next_k <= k_const(iteration+1);               end if;5��    M                     &      g               5�_�  ,  .          -  M       ����                                                                                                                                                                                                                                                                                                                i          N         N   "       V   '    f�     �  L  M                      -- Update kpw5��    L                     �%                     5�_�  -  /          .  M       ����                                                                                                                                                                                                                                                                                                                i          M         M   "       V   '    f�     �  M  O  f    �  M  N  f    5��    M                     &                     5�_�  .  0          /  N       ����                                                                                                                                                                                                                                                                                                                i          M         M   "       V   '    f�     �  M  O  g                  -- Update kpw5��    M                    &                     5�_�  /  =          0  N       ����                                                                                                                                                                                                                                                                                                                i          M         M   "       V   '    f�     �  M  O  g    5��    M                     &              	       �    M                     &                     5�_�  0  >  1      =  O        ����                                                                                                                                                                                                                                                                                                                i          Q          O           V        f�     �  N  O                  -- Update kpw   (        current_k <= k_const(iteration);   +        current_w <= w_vec(511 downto 480);5��    N                     &      k               5�_�  =  ?          >  M        ����                                                                                                                                                                                                                                                                                                                i          O          O           V        f�     �  L  P  e    �  M  N  e    5��    L                     �%              k       5�_�  >  @          ?  M       ����                                                                                                                                                                                                                                                                                                                i          @         S          V   "    f�   � �  M  P  h      (        current_k <= k_const(iteration);   +        current_w <= w_vec(511 downto 480);�  L  N  h              -- Update kpw5��    L                    &                     �    M                    &                     �    N                    K&                     5�_�  ?  A          @  N       ����                                                                                                                                                                                                                                                                                                                i          M         O                 f�3   � �  M  O  h      ,            current_k <= k_const(iteration);5��    M         	          "&      	              �    M                    $&                     �    M                    #&                     �    M                   "&                    �    M                   "&                    �    M                   "&                    5�_�  @  B          A  C       ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f�.     �  C  E  h    5��    C                     %%                     �    C                     %%                     5�_�  A  C          B  D        ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f�7     �  C  D           5��    C                     %%                     5�_�  B  D          C  G       ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f�:     �  G  I  i                  �  G  I  h    5��    G                     �%                     �    G                    �%                     �    G                    �%                     �    G                    �%                     �    G                   �%                    �    G                   �%                    �    G                   �%                    �    G                   �%                    �    G                   �%                    �    G                   �%                    5�_�  C  E          D  H       ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f�F     �  G  I  i                  next_k <= k_const5��    G                    �%                     5�_�  D  F          E  H       ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f�J     �  G  I  i                  next_k <= k_const()5��    G                    �%                     5�_�  E  G          F  H        ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f�L     �  G  I  i                   next_k <= k_const(1)5��    G                     �%                     5�_�  F  H          G  O   '    ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f�W     �  N  P  i      )            next_k <= k_const(iteration);5��    N  '                  _&                     5�_�  G  I          H  O   (    ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f�Z     �  N  P  j                  �  N  P  i    5��    N                     8&                     �    N                    D&                     �    N                   E&                    �    N                    H&                     �    N                	   G&             	       �    N         	          G&      	              �    N                   G&                    �    N                   R&                    5�_�  H  J          I  O       ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f�q     �  N  Q  j                  if iteration <= 615��    N                    V&                     �    N  #                  [&                     �    N  #                 [&                     �    O                    \&                    �    O                     \&                     5�_�  I  K          J  Q       ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f�}     �  Q  S  l                  �  Q  S  k    5��    Q                     �&                     �    Q                    �&                     �    Q                    �&                    �    Q                    �&                     5�_�  J  L          K  R       ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f��     �  Q  S  l              end if;5��    Q                    �&                     5�_�  K  M          L  P        ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f��     �  O  P           5��    O                     \&                     5�_�  L  N          M  P       ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f��     �  O  Q  k      +            next_k <= k_const(iteration+2);5��    O                    h&                     5�_�  M  O          N  Q       ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f��   � �  Q  S  k    5��    Q                     �&                     �    Q                     �&                     5�_�  N  P          O  K       ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f�     �  K  M  m                      �  K  M  l    5��    K                     	&                     �    K                    &                     �    K                    &                     �    K                    &                     �    K                   &                    �    K                   &                    �    K                
   &             
       5�_�  O  Q          P  L       ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f�     �  K  M  m                      enable <= 5��    K                    #&                     5�_�  P  R          Q  L       ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f�     �  K  M  m                      enable <= ''5��    K                    $&                     5�_�  Q  S          R  L       ����                                                                                                                                                                                                                                                                                                                i           �         =          v       f�    � �  K  M  m                      enable <= '0'5��    K                    &&                     5�_�  R  T          S  I       ����                                                                                                                                                                                                                                                                                                                i          0         7          v       f��     �  I  K  n                  �  I  K  m    5��    I                     �%              	       �    I                    �%                    �    I                	   �%             	       �    I                   �%                    5�_�  S  U          T  J       ����                                                                                                                                                                                                                                                                                                                i          0         7          v       f��     �  I  K  n                  enable <= 5��    I                    �%                     5�_�  T  V          U  J       ����                                                                                                                                                                                                                                                                                                                i          0         7          v       f��     �  I  K  n                  enable <= ''5��    I                    �%                     �    I                   �%                    5�_�  U  W          V  J       ����                                                                                                                                                                                                                                                                                                                i          0         7          v       f��     �  I  K  n                  enable <= '1'5��    I                    �%                     5�_�  V  X          W  B       ����                                                                                                                                                                                                                                                                                                                i          D         B          V       f��     �  A  B                  if rst = '0' then               enable <= '1';           end if;5��    A                     �$      E               5�_�  W  Y          X  G       ����                                                                                                                                                                                                                                                                                                                i          B         B          V       f�     �  G  J  l                  �  G  I  k    5��    G                     �%                     �    G                    �%                     �    G                    �%                     �    G                    �%                     �    G                	   �%             	       �    G         	          �%      	              �    G                   �%                    �    G                   �%                    �    G                   �%                    �    G                   �%                    �    G                   �%                     �    H                    �%                    �    H                     �%                     5�_�  X  Z          Y  H       ����                                                                                                                                                                                                                                                                                                                i          B         B          V       f�     �  G  I  m                  if iteration then5��    G                    �%                     �    G                   �%                    5�_�  Y  [          Z  L       ����                                                                                                                                                                                                                                                                                                                i          B         B          V       f�      �  K  L                          enable <= '0';5��    K                     &                     5�_�  Z  \          [  I        ����                                                                                                                                                                                                                                                                                                                i          B         B          V       f�"     �  H  J  l    �  I  J  l    5��    H                     �%                     5�_�  [  ]          \  J        ����                                                                                                                                                                                                                                                                                                                i          B         B          V       f�#   � �  I  K  m       5��    I                     �%                     �    I                    �%                    �    I                    �%                     5�_�  \  ^          ]  L       ����                                                                                                                                                                                                                                                                                                                i          H         J          V       f�~     �  K  M  n                      �  K  M  m    5��    K                     &                     �    K                    (&                     �    K                    *&                     �    K                    )&                     �    K                   (&                    �    K                   (&                    �    K                
   (&             
       5�_�  ]  _          ^  L       ����                                                                                                                                                                                                                                                                                                                i          H         J          V       f�     �  K  M  n                      enable <= 5��    K                    2&                     5�_�  ^  `          _  L       ����                                                                                                                                                                                                                                                                                                                i          H         J          V       f�     �  K  M  n                      enable <= ''5��    K                    3&                     5�_�  _  f          `  L       ����                                                                                                                                                                                                                                                                                                                i          H         J          V       f�   � �  K  M  n                      enable <= '0'5��    K                    5&                     5�_�  `  g  a      f  R   ,    ����                                                                                                                                                                                                                                                                                                                i          H         J          V       f�M     �  Q  S  n      /                next_k <= k_const(iteration+2);5��    Q  ,                 �&                    5�_�  f  h          g  Q       ����                                                                                                                                                                                                                                                                                                                i          H         J          V       f�P   � �  P  R  n      #            if iteration <= 61 then5��    P                   �&                    5�_�  g  i          h  E       ����                                                                                                                                                                                                                                                                                                                i          H         J          V       f��   � �  D  E          !            next_k <= k_const(1);5��    D                     >%      "               5�_�  h  j          i         ����                                                                                                                                                                                                                                                                                                                i          J         K          v       f�_     �      m      L    get_k: reg32 port map (rst, clk, enable, k_const(0), next_k, current_k);5��                        �      M       P       5�_�  i  k          j  P       ����                                                                                                                                                                                                                                                                                                                i          R         O          V       f�     �  N  P  j                  -- Update kpw�  O  P          #            if iteration <= 62 then   /                next_k <= k_const(iteration+1);               end if;5��    O                     d&      h               �    N                   V&                    �    N                    X&                     �    N                    W&                     �    N                	   V&             	       �    N         	          V&      	              �    N                   V&                    �    N                    e&                     �    N                    d&                     �    N                   c&                    �    N                   c&                    �    N                   c&                    5�_�  j  l          k  O        ����                                                                                                                                                                                                                                                                                                                i          P         O          V       f�     �  N  P  j                   current_k <= k_const5��    N                     j&                     5�_�  k  m          l  O   !    ����                                                                                                                                                                                                                                                                                                                i          P         O          V       f�     �  N  P  j      "            current_k <= k_const()5��    N  !                  k&                     �    N  !              	   k&             	       �    N  !       	          k&      	              �    N  !              	   k&             	       5�_�  l  n          m  O   +    ����                                                                                                                                                                                                                                                                                                                i          P         O          V       f�   � �  N  P  j      +            current_k <= k_const(iteration)5��    N  +                  u&                     5�_�  m  o          n  O       ����                                                                                                                                                                                                                                                                                                                i          P         O          V       f�     �  N  O          ,            current_k <= k_const(iteration);5��    N                     J&      -               5�_�  n  p          o  Q        ����                                                                                                                                                                                                                                                                                                                i          O         O          V       f�   � �  Q  S  i    �  Q  R  i    5��    Q                     �&              -       5�_�  o  q          p  P       ����                                                                                                                                                                                                                                                                                                                i          O         O          V       f�     �  O  P          /            current_w <= w_vec(511 downto 480);5��    O                     K&      0               5�_�  p  r          q  Q       ����                                                                                                                                                                                                                                                                                                                i          O         O          V       f�   � �  Q  S  i    �  Q  R  i    5��    Q                     �&              0       5�_�  q  s          r  R       ����                                                                                                                                                                                                                                                                                                                i          O         O          V       f��     �  Q  R          /            current_w <= w_vec(511 downto 480);5��    Q                     �&      0               5�_�  r  t          s  P        ����                                                                                                                                                                                                                                                                                                                i          O         O          V       f��   � �  O  Q  i    �  P  Q  i    5��    O                     K&              0       5�_�  s  u          t   �       ����                                                                                                                                                                                                                                                                                                                i             6       �          v   >    f��     �   �   �  j      #    signal iteration: integer := 0;5��    �                     �                     �    �   $                 �                    �    �   %                 �                    �    �   &                 �                    �    �   '                 �                    5�_�  t  v          u   �   $    ����                                                                                                                                                                                                                                                                                                                i             6       �          v   >    f��     �   �   �  j      )    signal iteration: integer range  to ;5��    �   $                  �                     5�_�  u  w          v   �   )    ����                                                                                                                                                                                                                                                                                                                i             6       �          v   >    f��   � �   �   �  j      *    signal iteration: integer range 0 to ;5��    �   )                  �                     5�_�  v  x          w   T       ����                                                                                                                                                                                                                                                                                                                i             6       �          v   >    f�3     �   S   U  j      !    count <= to_integer(counter);5��    S          
           	      
               5�_�  w  y          x   T       ����                                                                                                                                                                                                                                                                                                                i             6       �          v   >    f�4     �   S   U  j          count <= (counter);5��    S                     	                     5�_�  x  z          y   T       ����                                                                                                                                                                                                                                                                                                                i             6       �          v   >    f�7     �   S   U  j          count <= counter);5��    S                                          5�_�  y  {          z   B       ����                                                                                                                                                                                                                                                                                                                i             6       �          v   >    f�?     �   A   C  j      B        count : out integer       -- 6-bit count output (64 steps)5��    A                    i                    �    A                     l                     �    A                     k                     �    A                     j                     �    A                    i                    �    A                    i                    �    A                    i                    5�_�  z  |          {   B       ����                                                                                                                                                                                                                                                                                                                i             6       �          v   >    f�B     �   A   C  j      C        count : out unsigned       -- 6-bit count output (64 steps)5��    A                     q                     5�_�  {  }          |   B       ����                                                                                                                                                                                                                                                                                                                i             6       �          v   >    f�E     �   A   C  j      E        count : out unsigned()       -- 6-bit count output (64 steps)5��    A                     r                     �    A                     t                     �    A                     s                     �    A                    r                    �    A                    t                    �    A                    t                    �    A                    t                    5�_�  |  ~          }   �       ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f�j     �   �   �  j      ,    signal iteration: integer range 0 to 63;5��    �                    �                    �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�  }            ~   �       ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f�l     �   �   �  j          signal iteration: unsigned;5��    �                     �                     5�_�  ~  �             �       ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f�n     �   �   �  j      !    signal iteration: unsigned();5��    �                     �                     �    �   !                 �                    �    �   !                 �                    �    �   !                 �                    5�_�    �          �   �       ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f�     �   �   �  j      F            count : out integer       -- 6-bit count output (64 steps)5��    �                    �                    �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f�     �   �   �  j      G            count : out unsigned       -- 6-bit count output (64 steps)5��    �                      �                     5�_�  �  �          �   �   !    ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f�     �   �   �  j      I            count : out unsigned()       -- 6-bit count output (64 steps)5��    �   !                  �                     �    �   #                 �                    �    �   #                 �                    �    �   #                 �                    5�_�  �  �          �  G       ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f�     �  F  H  j      "            if iteration = 62 then5��    F                    �%                     5�_�  �  �          �  G       ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f�     �  F  H  j      #            if (iteration = 62 then5��    F                    �%      $       %       5�_�  �  �          �  G       ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f�     �  F  H  j      $            if (iteration) = 62 then5��    F                    �%                     �    F                   �%                    5�_�  �  �          �  J       ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f�     �  I  K  j      "            if iteration = 63 then5��    I                    &                     5�_�  �  �          �  J       ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f�     �  I  K  j      #            if (iteration = 63 then5��    I                    �%      $       %       5�_�  �  �          �  J       ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f�     �  I  K  j      $            if (iteration) = 63 then5��    I                    &                     �    I                    &                     �    I                
   &             
       �    I         
          &      
              �    I                
   &             
       5�_�  �  �          �  R   !    ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f�     �  Q  S  j      ,            current_k <= k_const(iteration);5��    Q  !                  �&                     �    Q  "                  �&                     �    Q  !              
   �&             
       �    Q  !       
          �&      
              �    Q  !                 �&                    5�_�  �  �          �  R   ,    ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f�   � �  Q  S  j      7            current_k <= k_const(to_integer(iteration);5��    Q                    �&      8       9       5�_�  �  �  �      �     6    ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f��     �              O    -- get_k: reg32 port map (rst, clk, enable, k_const(0), next_k, current_k);5��                               P               5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f��     �               5��                                              5�_�  �  �          �  N       ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f��     �  M  N          /            current_w <= w_vec(511 downto 480);5��    M                     (&      0               5�_�  �  �          �  N       ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f��   � �  N  P  g    �  N  O  g    5��    N                     8&              0       5�_�  �  �          �  !   %    ����                                                                                                                                                                                                                                                                                                                i          !   %      (   (          (    f��   � �     "  h      :    get_aout: adder32 port map (h0, a, haso(31 downto 0));�     )  h      >    get_aout: adder32 port map (h0, a_reg, haso(31 downto 0));   ?    get_bout: adder32 port map (h1, b_reg, haso(63 downto 32));   ?    get_cout: adder32 port map (h2, c_reg, haso(95 downto 64));   @    get_dout: adder32 port map (h3, d_reg, haso(127 downto 96));   A    get_eout: adder32 port map (h4, e_reg, haso(159 downto 128));   A    get_fout: adder32 port map (h5, f_reg, haso(191 downto 160));   A    get_gout: adder32 port map (h6, g_reg, haso(223 downto 192));   A    get_hout: adder32 port map (hv, h_reg, haso(255 downto 224));5��       %                  <!                     �    !  %                  w!                     �    "  %                  �!                     �    #  %                  �!                     �    $  %                  ,"                     �    %  %                  j"                     �    &  %                  �"                     �    '  %                  �"                     �       %                  <!                     �    !  %                  x!                     �    "  %                  �!                     �    #  %                  �!                     �    $  %                  0"                     �    %  %                  o"                     �    &  %                  �"                     �    '  %                  �"                     5�_�  �  �  �      �   �       ����                                                                                                                                                                                                                                                                                                                i          !   %      (   (          (    f��     �   �   �          +    signal next_k: bit_vector(31 downto 0);5��    �                      )      ,               5�_�  �  �  �      �   A       ����                                                                                                                                                                                                                                                                                                                i              %      '   (          (    f      �   @   B  g      K        clk, rst, enable: in bit;                            -- Clock input5��    @                                          5�_�  �  �          �   B       ����                                                                                                                                                                                                                                                                                                                i              %      '   (          (    f      �   A   C  h          �   A   C  g    5��    A                      M              	       �    A                     M                    �    A                    X                    �    A                    Y                    �    A                    Y                    �    A                    [                    �    A                    b                    5�_�  �  �          �   O       ����                                                                                                                                                                                                                                                                                                                j          !   %      (   (          (    f U     �   O   Q  i                  �   O   Q  h    5��    O                      �                     �    O                  	   �              	       �    O                     �                     5�_�  �  �          �   P       ����                                                                                                                                                                                                                                                                                                                k          "   %      )   (          (    f Z     �   O   Q  i                  done <= 5��    O                     �                     5�_�  �  �          �   P       ����                                                                                                                                                                                                                                                                                                                k          "   %      )   (          (    f Z     �   O   Q  i                  done <= ''5��    O                     �                     �    O                    �                    5�_�  �  �          �   P       ����                                                                                                                                                                                                                                                                                                                k          "   %      )   (          (    f \     �   O   Q  i                  done <= '0'5��    O                     �                     5�_�  �  �          �   Q       ����                                                                                                                                                                                                                                                                                                                k          "   %      )   (          (    f d     �   P   R  i      4        elsif rising_edge(clk) and enable = '1' then5��    P                     �                     5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                k          "   %      )   (          (    f p     �   Q   S  j                  �   Q   S  i    5��    Q                      �                     �    Q                     �                     5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                l          #   %      *   (          (    f z     �   Q   S  j                  if counter = 5��    Q                     �                     5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                l          #   %      *   (          (    f {     �   Q   S  j                  if counter = ""5��    Q                     �                     5�_�  �  �          �   R   !    ����                                                                                                                                                                                                                                                                                                                l          #   %      *   (          (    f      �   Q   S  j      !            if counter = "000000"5��    Q   !                  �                     �    Q   %                  �                     �    Q   $                  �                     �    Q   #                  �                     �    Q   "                  �                     �    Q   !                  �                     �    Q                     �                     �    Q                     �                     5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                l          #   %      *   (          (    f �     �   Q   S  j                  if counter = 5��    Q                     �                     5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                l          #   %      *   (          (    f �     �   Q   S  j                  if counter = ()5��    Q                     �                     �    Q                    �                    �    Q                    �                    �    Q                    �                    �    Q                    �                    5�_�  �  �          �   R   (    ����                                                                                                                                                                                                                                                                                                                l          #   %      *   (          (    f �     �   Q   T  j      (            if counter = (others => '0')5��    Q   (                  �                     �    Q   -                  �                     �    Q   -                 �                     �    R                     �                    �    R                      �                     5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                m          $   %      +   (          (    f �     �   Q   S  k      -            if counter = (others => '0') then5��    Q                     �                     �    Q                     �                     �    Q                    �                    �    Q                     �                     �    Q                 
   �             
       �    Q          
          �      
              �    Q                 
   �             
       5�_�  �  �          �   R   #    ����                                                                                                                                                                                                                                                                                                                m          $   %      +   (          (    f �     �   Q   S  k      (            if counter = to_integer then5��    Q   #                  �                     5�_�  �  �          �   R   $    ����                                                                                                                                                                                                                                                                                                                m          $   %      +   (          (    f �     �   Q   S  k      *            if counter = to_integer() then5��    Q   #                  �                     �    Q          	           �      	               �    Q                     �                     �    Q                    �                    �    Q                     �                     �    Q                    �                    �    Q                    �                    �    Q                    �                    5�_�  �  �          �   R   !    ����                                                                                                                                                                                                                                                                                                                m          $   %      +   (          (    f �     �   Q   S  k      &            if counter = unsigned then5��    Q   !                  �                     5�_�  �  �          �   R   "    ����                                                                                                                                                                                                                                                                                                                m          $   %      +   (          (    f �     �   Q   S  k      (            if counter = unsigned() then5��    Q   "                  �                     5�_�  �  �          �   S        ����                                                                                                                                                                                                                                                                                                                m          $   %      +   (          (    f �     �   R   T  k       5��    R                      �                     �    R                                          �    R                                        5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                m          $   %      +   (          (    f �     �   R   T  k                      done <= 5��    R                                          5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                m          $   %      +   (          (    f �     �   R   T  k                      done <= ''5��    R                                          5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                m          $   %      +   (          (    f �     �   R   T  k                      done <= '0'5��    R                                          5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                m          $   %      +   (          (    f �     �   R   T  k                      done <= '0';5��    R                                        5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                m          $   %      +   (          (    f �     �   R   U  k                      done <= '1';5��    R                                         �    S                    %                    5�_�  �  �          �   U       ����                                                                                                                                                                                                                                                                                                                n          %   %      ,   (          (    f �     �   T   V  l      #            counter <= counter + 1;5��    T                     6                     �    T                    6                    5�_�  �  �          �   U       ����                                                                                                                                                                                                                                                                                                                n          %   %      ,   (          (    f �     �   U   W  m                      �   U   W  l    5��    U                      R                     �    U                     b                     �    U                     R                    �    U                     b                     �    U                    d                    5�_�  �  �  �      �   R       ����                                                                                                                                                                                                                                                                                                                o          &   %      -   (          (    f �     �   Q   S  m      *            if counter = unsigned(63) then5��    Q                     �                     5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                o          &   %      -   (          (    f �     �   Q   S  m      "            if counter = (63) then5��    Q                     �                     5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                o          &   %      -   (          (    f �     �   Q   S  m      !            if counter = 63) then5��    Q                     �                     5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                o          &   %      -   (          (    f �     �   Q   S  m                   if counter = 63 then5��    Q                     �                     5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                o          &   %      -   (          (    f �     �   Q   S  m      !            if (counter = 63 then5��    Q                     �      "       #       5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                o          &   %      -   (          (    f �     �   Q   S  m      "            if (counter) = 63 then5��    Q                     �                     �    Q                     �                     �    Q                 
   �             
       �    Q          
          �      
              �    Q                 
   �             
       5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                o          &   %      -   (          (    f �     �   S   U  n                      �   S   U  m    5��    S                                           �    S                     +                     �    S                     .                     �    S                     -                     �    S                     ,                     �    S                    +                    �    S                    +                    �    S                    +                    5�_�  �  �          �   T       ����                                                                                                                                                                                                                                                                                                                p          '   %      .   (          (    f �   � �   S   T                          counter5��    S                                           5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                o          &   %      -   (          (    f     �   �   �  m      "    signal enable: bit := not rst;5��    �                    C                    5�_�  �  �  �      �   �       ����                                                                                                                                                                                                                                                                                                                o           �          �          v       f%     �   �   �  m      !    signal ended: bit := not rst;5��    �                     M                     5�_�  �  �          �     ,    ����                                                                                                                                                                                                                                                                                                                o           �          �          v       f9     �      m      I    shf_w: shift_reg512 port map (rst, clk, enable, next_w, msgi, w_vec);5��      ,              	   �             	       5�_�  �  �          �     .    ����                                                                                                                                                                                                                                                                                                                o           �          �          v       f?     �      m      A    counter: counter_6bit port map (clk, rst, enable, iteration);5��      .                 F                    �      .                  F                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                o           �          �          v       fH     �   �   �  m      O            clk, rst, enable: in bit;                            -- Clock input5��    �                     �                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                o           �          �          v       fI     �   �   �  m      N            clk, rst enable: in bit;                            -- Clock input5��    �                     �                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                o           �          �          v       fI     �   �   �  m      M            clk, rstenable: in bit;                            -- Clock input5��    �                     �                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                o           �          �          v       fK     �   �   �  n              �   �   �  m    5��    �                      3                     �    �                     3                    5�_�  �  �          �     .    ����                                                                                                                                                                                                                                                                                                                o           �          �          v       fk     �      n      ;    counter: counter_6bit port map (clk, rst, , iteration);5��      .                  Y                     �      0                 [                    5�_�  �  �          �     *    ����                                                                                                                                                                                                                                                                                                                o             *      %   /          /    fy     �      n      ;    a_register: reg32 port map (rst, clk, , h0, av, a_reg);�    &  n      A    a_register: reg32 port map (rst, clk, enable, h0, av, a_reg);   A    b_register: reg32 port map (rst, clk, enable, h1, bv, b_reg);   A    c_register: reg32 port map (rst, clk, enable, h2, cv, c_reg);   A    d_register: reg32 port map (rst, clk, enable, h3, dv, d_reg);   A    e_register: reg32 port map (rst, clk, enable, h4, ev, e_reg);   A    f_register: reg32 port map (rst, clk, enable, h5, fv, f_reg);   A    g_register: reg32 port map (rst, clk, enable, h6, gv, g_reg);   A    h_register: reg32 port map (rst, clk, enable, h7, hv, h_reg);5��      *                  �                     �      *                  �                     �      *                                        �       *                  K                      �    !  *                  �                      �    "  *                  �                      �    #  *                  �                      �    $  *                  ;!                     �      *               	   �              	       �      *               	   �              	       �      *               	   !               	       �       *               	   f               	       �    !  *               	   �               	       �    "  *               	   �               	       �    #  *               	   5!              	       �    $  *               	   z!              	       5�_�  �  �          �  H       ����                                                                                                                                                                                                                                                                                                                o             *      %   /          /    f�     �  G  H                      enable <= '0';5��    G                     R%                     5�_�  �  �          �  I       ����                                                                                                                                                                                                                                                                                                                o             *      %   /          /    f�     �  H  I                      enable <= '1';5��    H                     v%                     5�_�  �  �          �  J       ����                                                                                                                                                                                                                                                                                                                o             *      %   /          /    f�     �  I  J                          enable <= '0';5��    I                     �%                     5�_�  �  �          �  L       ����                                                                                                                                                                                                                                                                                                                o             *      %   /          /    f�     �  K  L                          enable <= '0';5��    K                     �%                     5�_�  �  �          �  Q       ����                                                                                                                                                                                                                                                                                                                o             *      %   /          /    f�     �  P  R  j      /            current_w <= w_vec(511 downto 480);5��    P                    3&                     5�_�  �  �          �  R       ����                                                                                                                                                                                                                                                                                                                o             *      %   /          /    f�     �  Q  S  j      8            current_k <= k_const(to_integer(iteration));5��    Q                    _&                     5�_�  �  �          �  Q       ����                                                                                                                                                                                                                                                                                                                o             *      %   /          /    f�     �  P  S  k              �  P  R  j    5��    P                     +&              	       �    P                     +&                     �    P                    +&              	       �    Q                    4&                     5�_�  �  �          �  V        ����                                                                                                                                                                                                                                                                                                                o          D         P          V       f�     �  U  V                  end process;5��    U                     �&                     5�_�  �  �          �  U        ����                                                                                                                                                                                                                                                                                                                o          D         P          V       f�     �  T  U           5��    T                     �&                     5�_�  �  �          �  D       ����                                                                                                                                                                                                                                                                                                                o          P         D          V       f�     �  C  D              process(clk, rst)   	    begin           if rst = '1' then               done <= '0';   #        elsif rising_edge(clk) then   .            if to_integer(iteration) = 62 then               end if;   .            if to_integer(iteration) = 63 then                   done <= '1';               end if;                   end if;5��    C                     �$      ,              5�_�  �  �          �  D        ����                                                                                                                                                                                                                                                                                                                o          D         D          V       f�     �  C  D           5��    C                     �$                     5�_�  �  �          �  D       ����                                                                                                                                                                                                                                                                                                                o          D         F                 f�     �  C  E  [              done <= ended;5��    C                    %                     5�_�  �  �          �  E       ����                                                                                                                                                                                                                                                                                                                o          D         F                 f�     �  D  F  [      +        current_w <= w_vec(511 downto 480);5��    D                    %                     5�_�  �  �          �  F       ����                                                                                                                                                                                                                                                                                                                o          D         F                 f�   � �  E  G  [      4        current_k <= k_const(to_integer(iteration));5��    E                    >%                     5�_�  �  �  �      �  '   %    ����                                                                                                                                                                                                                                                                                                                o          '   %      .   %          %    f�"   � �  &  (  [      :    get_aout: adder32 port map (h0, a, haso(31 downto 0));�  &  /  [      ;    get_aout: adder32 port map (h0, av, haso(31 downto 0));   <    get_bout: adder32 port map (h1, bv, haso(63 downto 32));   <    get_cout: adder32 port map (h2, cv, haso(95 downto 64));   =    get_dout: adder32 port map (h3, dv, haso(127 downto 96));   >    get_eout: adder32 port map (h4, ev, haso(159 downto 128));   >    get_fout: adder32 port map (h5, fv, haso(191 downto 160));   >    get_gout: adder32 port map (h6, gv, haso(223 downto 192));   >    get_hout: adder32 port map (hv, hv, haso(255 downto 224));5��    &  %                  �!                     �    '  %                  �!                     �    (  %                  2"                     �    )  %                  n"                     �    *  %                  �"                     �    +  %                  �"                     �    ,  %                  '#                     �    -  %                  e#                     �    &  %                  �!                     �    '  %                  �!                     �    (  %                  :"                     �    )  %                  z"                     �    *  %                  �"                     �    +  %                  �"                     �    ,  %                  ?#                     �    -  %                  �#                     5�_�  �  �  �      �   R   &    ����                                                                                                                                                                                                                                                                                                                o           R   (       T          V   (    f�   � �   Q   S  [      ,            if to_integer(counter) = 63 then5��    Q   &                 �                    5�_�  �  �          �   X       ����                                                                                                                                                                                                                                                                                                                o           R   (       T          V   (    fR     �   Z   ]  ^              �   Y   \  ]          if�   X   [  \          �   X   Z  [    5��    X                      �                     �    X                      �                     �    X                     �                     �    Y                     �                     �    Y                    �                    �    Y                    �                    �    Y                    �                    �    Y                    �                    �    Y                    �                    �    Y                    �                     �    Z                      �                      �    Z                    �                     5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                s           Z          Z          v       fW     �   Y   [  _          if condition then5��    Y          	          �      	              5�_�  �  �          �   [        ����                                                                                                                                                                                                                                                                                                                s           Z          \          V       f[     �   [   ]  _          end generate �   Z   ]  ^              �   Y   \  ]          if rs then�   Z   [                         end if;5��    Z                      �                     �    Y          
          �      
              �    Y                     �                     �    Y                    �                    �    Y                    �                    �    Y                    �                    �    Y                    �                    �    Y                     �                     �    Z                      �                      �    Z                    �                     �    [                     �                     5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                s           Z          Z          v       f`     �   Z   [  _    �   [   ]  _           end generate generate_label;�   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Z   [  _    �   Y   [  _      )    generate_label: if condition generate5��    Y                    �                    �    [                    �                    �    Y                     �                     �    [                    �                    �    Y                     �                     �    [                    �                    �    Y                     �                     �    [                    �                    �    Y                     �                     �    [                    �                    �    Y                     �                     �    [                    �                    �    Y                     �                     �    [                    �                    �    Y                     �                     �    [                    �                    �    Y                     �                     �    [                    �                    �    Y                     �                     �    [                     �                     �    Y                     �                     �    [                     �                     �    Y                     �                     �    [                    �                    �    Y                     �                     �    [                    �                    �    Y                     �                     �    [                    �                    �    Y                     �                     �    [                    �                    �    Y   	                  �                     �    [                    �                    �    Y   
                  �                     �    [                    �                    �    Y                     �                     �    [                    �                    �    Y                     �                     �    [                 	   �             	       �    Y                     �                     �    [          	       
   �      	       
       5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                s           Z          Z          v       fm     �   Y   [  _      %    done_check: if condition generate5��    Y          	          �      	              �    Y                     �                     �    Y                    �                    �    Y                    �                    �    Y                    �                    5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                s           Z          Z          v       fp     �   Y   [  _      "    done_check: if rst =  generate5��    Y                     �                     5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                s           Z          Z          v       fq     �   Y   [  _      $    done_check: if rst = '' generate5��    Y                     �                     5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                s           Z          Z          v       fr     �   Y   [  _      %    done_check: if rst = '0' generate5��    Y                     �                     �    Y   "                  �                     �    Y   !              
   �             
       �    Y   !       
          �      
              �    Y   !              
   �             
       5�_�  �  �          �   Z   +    ����                                                                                                                                                                                                                                                                                                                s           Z          Z          v       fv     �   Y   [  _      4    done_check: if rst = '0' and to_integer generate5��    Y   +                  �                     5�_�  �  �          �   Z   ,    ����                                                                                                                                                                                                                                                                                                                s           Z          Z          v       fv     �   Y   [  _      6    done_check: if rst = '0' and to_integer() generate5��    Y   ,                  �                     �    Y   -                  �                     �    Y   ,                 �                    �    Y   /                  �                     �    Y   .                  �                     �    Y   -                  �                     �    Y   ,                 �                    �    Y   2                  �                     �    Y   1                  �                     �    Y   0                  �                     �    Y   /                  �                     �    Y   .                  �                     �    Y   -                  �                     �    Y   ,                 �                    �    Y   ,                 �                    �    Y   ,                 �                    5�_�  �  �          �   Z   4    ����                                                                                                                                                                                                                                                                                                                s           Z          Z          v       fy     �   Y   [  _      =    done_check: if rst = '0' and to_integer(counter) generate5��    Y   4                  �                     5�_�  �  �          �   Z   8    ����                                                                                                                                                                                                                                                                                                                s           Z          Z          v       f�     �   Y   [  _      B    done_check: if rst = '0' and to_integer(counter) = 62 generate5��    Y   8                 �                    5�_�  �  �          �   [       ����                                                                                                                                                                                                                                                                                                                s           Z          Z          v       f�     �   Z   \  _              5��    Z                     �                     �    Z   
                  �                     �    Z   	                  �                     �    Z                 
   �             
       �    Z                     �                     �    Z                     �                     �    Z                     �                     �    Z                     �                     �    Z                     �                     �    Z                     �                     �    Z                     �                     �    Z   
                  �                     �    Z   	                  �                     �    Z                    �                    �    Z                     �                     �    Z   
                  �                     �    Z   	                  �                     �    Z                    �                    �    Z                    �                    �    Z                    �                    �    Z                    �                    5�_�  �  �          �   [       ����                                                                                                                                                                                                                                                                                                                s           Z          Z          v       f�     �   Z   \  _              done <= 5��    Z                     �                     5�_�  �  �          �   [       ����                                                                                                                                                                                                                                                                                                                s           Z          Z          v       f�     �   Z   \  _              done <= ''5��    Z                     �                     5�_�  �  �          �   [       ����                                                                                                                                                                                                                                                                                                                s           Z          Z          v       f�     �   Z   \  _              done <= '1'5��    Z                     �                     5�_�  �  �          �   R        ����                                                                                                                                                                                                                                                                                                                s           R          T          V       f�     �   Q   R          ,            if to_integer(counter) = 62 then                   done <= '1';               else5��    Q                      �      [               5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                p           R          R          V       f�     �   R   S                      end if;5��    R                      �                     5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                o           R          R          V       f�   � �   Q   S  [      '                counter <= counter + 1;5��    Q                     �                     5�_�  �  �  �      �   V       ����                                                                                                                                                                                                                                                                                                                o           X          V          V       f     �   U   W  [      B    done_check: if rst = '0' and to_integer(counter) = 63 generate5��    U                     $                     5�_�  �  �          �   X       ����                                                                                                                                                                                                                                                                                                                o           X          V          V       fO     �   W   Y  [          end generate done_check;5��    W                    t                    5�_�  �            �   V   .    ����                                                                                                                                                                                                                                                                                                                o           X          V          V       fV     �   U   W  [      6    if rst = '0' and to_integer(counter) = 63 generate5��    U   .                 N                    5�_�  �    �         P       ����                                                                                                                                                                                                                                                                                                                o           X   
       V          V       f�     �   P   R  \              elsif�   O   R  [                  done <= '0';5��    O                    �                     �    P                    �                    �    P   	                  �                     �    P                    �                    �    P   
                  �                     �    P   	                  �                     �    P                    �                    �    P                    �                    �    P                    �                    �    P                     �                     �    P                 
   �             
       �    P          
          �      
              �    P                 
   �             
       5�_�                 Q       ����                                                                                                                                                                                                                                                                                                                p           Y   
       W          V       f�     �   P   R  \              elsif to_integer5��    P                     �                     5�_�                 Q       ����                                                                                                                                                                                                                                                                                                                p           Y   
       W          V       f�     �   P   R  \              elsif to_integer()5��    P                     �                     �    P                    �                    �    P                    �                    �    P                    �                    5�_�                 Q   !    ����                                                                                                                                                                                                                                                                                                                p           Y   
       W          V       f�     �   P   R  \      !        elsif to_integer(counter)5��    P   !                  �                     �    P   "                 �                    5�_�                 Q   &    ����                                                                                                                                                                                                                                                                                                                p           Y   
       W          V       f�     �   Q   S  ]                  done�   P   S  \      &        elsif to_integer(counter) = 635��    P   &                  �                     �    P   +                  �                     �    P   +                 �              	       �    Q                     �                    �    Q                     �                     �    Q                     �                     �    Q                    �                    �    Q                    �                    �    Q                    �                    �    Q                     �                     �    Q                    �                    5�_�                 R       ����                                                                                                                                                                                                                                                                                                                q           Z   
       X          V       f     �   Q   S  ]                  done <= 1;5��    Q                     �                     5�_�                 R       ����                                                                                                                                                                                                                                                                                                                q           Z   
       X          V       f     �   Q   S  ]                  done <= ;5��    Q                     �                     5�_�    	             R       ����                                                                                                                                                                                                                                                                                                                q           Z   
       X          V       f     �   Q   S  ]                  done <= '';5��    Q                     �                     5�_�    
          	   X        ����                                                                                                                                                                                                                                                                                                                q           Z   
       X          V       f   � �   W   X          2    if rst = '0' and to_integer(counter) = 63 then           done <= '1';       end if;    5��    W                      e      U               5�_�  	            
  %   %    ����                                                                                                                                                                                                                                                                                                                m          %   %      ,   (          (    f`   � �  $  &  Y      :    get_aout: adder32 port map (h0, a, haso(31 downto 0));�  $  -  Y      >    get_aout: adder32 port map (h0, a_reg, haso(31 downto 0));   ?    get_bout: adder32 port map (h1, b_reg, haso(63 downto 32));   ?    get_cout: adder32 port map (h2, c_reg, haso(95 downto 64));   @    get_dout: adder32 port map (h3, d_reg, haso(127 downto 96));   A    get_eout: adder32 port map (h4, e_reg, haso(159 downto 128));   A    get_fout: adder32 port map (h5, f_reg, haso(191 downto 160));   A    get_gout: adder32 port map (h6, g_reg, haso(223 downto 192));   A    get_hout: adder32 port map (hv, h_reg, haso(255 downto 224));5��    $  %                  �!                     �    %  %                  �!                     �    &  %                  "                     �    '  %                  @"                     �    (  %                  }"                     �    )  %                  �"                     �    *  %                  �"                     �    +  %                  7#                     �    $  %                  �!                     �    %  %                  �!                     �    &  %                  "                     �    '  %                  C"                     �    (  %                  �"                     �    )  %                  �"                     �    *  %                  �"                     �    +  %                  >#                     5�_�  
  Z           2       ����                                                                                                                                                                                                                                                                                                                m           <          Z          V       f�   � �   1   3  Y                  vector <= d;5��    1                    �                    5�_�    [          Z   2       ����                                                                                                                                                                                                                                                                                                                m          %   %      ,   (          (    f(h�   � �   1   3  Y                  q <= d;5��    1                    �                    �    1                     �                     �    1                     �                     �    1                    �                    �    1                    �                    �    1                    �                    5�_�  Z  \          [   �       ����                                                                                                                                                                                                                                                                                                                M                                            f=�     �   �   �  [          signal haso0: bit_vector�   �   �  Z          �   �   �  Y    5��    �                                           �    �                                           �    �                                          �    �                                           �    �                     0                     �    �                     /                     �    �                    .                    �    �                     0                     �    �                     /                     �    �                 
   .             
       �    �                     7                     �    �                     6                     �    �                     5                     �    �                     4                     �    �                     3                     �    �                     2                     �    �                     1                     �    �                     0                     �    �                     /                     �    �                 
   .             
       �    �          
          .      
              �    �                 
   .             
       5�_�  [  ]          \   �       ����                                                                                                                                                                                                                                                                                                                M                                            f=     �   �   �  [          signal haso0: bit_vector5��    �                     8                     5�_�  \  ^          ]   �       ����                                                                                                                                                                                                                                                                                                                M                                            f=     �   �   �  [          signal haso0: bit_vector()5��    �                     9                     �    �                     <                    �    �                     <                    �    �                     <                    5�_�  ]  d          ^   �   )    ����                                                                                                                                                                                                                                                                                                                M                                            f=	     �   �   �  [      )    signal haso0: bit_vector(31 downto 0)5��    �   )                  E                     5�_�  ^  h  _      d   �   )    ����                                                                                                                                                                                                                                                                                                                M                                            f=     �   �   �  [    �   �   �  [    5��    �                      G              -      5�_�  d  i  g      h   �       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �   �   �  b      *    signal haso0: bit_vector(31 downto 0);5��    �                    V                    5�_�  h  j          i   �       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �   �   �  b      *    signal haso0: bit_vector(31 downto 0);5��    �                    �                    5�_�  i  k          j   �       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �   �   �  b      *    signal haso0: bit_vector(31 downto 0);5��    �                    �                    5�_�  j  l          k   �       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �   �   �  b      *    signal haso0: bit_vector(31 downto 0);5��    �                    �                    5�_�  k  m          l   �       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �   �   �  b      *    signal haso0: bit_vector(31 downto 0);5��    �                                        5�_�  l  n          m   �       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �   �   �  b      *    signal haso0: bit_vector(31 downto 0);5��    �                    -                    5�_�  m  o          n   �       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �   �   �  b      *    signal haso0: bit_vector(31 downto 0);5��    �                    X                    5�_�  n  q          o  5       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �  5  7  b    5��    5                     �$                     �    5                     �$                     5�_�  o  r  p      q  6        ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �  6  8  d          �  6  8  c    5��    6                     �$                     �    6                     �$                     5�_�  q  s          r  7       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �  6  8  d          haso0 <= haso5��    6                    �$                     5�_�  r  t          s  7       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �  6  8  d          haso0 <= haso()5��    6                    �$                     5�_�  s  u          t  7       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �  6  8  d          haso0 <= haso( downto )5��    6                    �$                     5�_�  t  v          u  7       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �  6  8  d          haso0 <= haso( downto );5��    6                    �$                     5�_�  u  x          v  7       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �  7  ?  d    �  7  8  d    5��    7                     �$              �       5�_�  v  y  w      x  8       ����                                                                                                                                                                                                                                                                                                                M          8         >                 f=�     �  7  ?  k          haso0 <= haso();       haso0 <= haso();       haso0 <= haso();       haso0 <= haso();       haso0 <= haso();       haso0 <= haso();       haso0 <= haso();5��    7                   �$                    �    8                   �$                    �    9                   �$                    �    :                   %                    �    ;                   #%                    �    <                   8%                    �    =                   M%                    5�_�  x  z          y  7       ����                                                                                                                                                                                                                                                                                                                M          .   -      5   8          8    f=     �  6  @  k   	       haso0 <= haso();       haso1 <= haso();       haso2 <= haso();       haso3 <= haso();       haso4 <= haso();       haso5 <= haso();       haso6 <= haso();       haso7 <= haso();    �  7  8  k    5��    6                    �$                     �    7                    �$                     �    8                    %                     �    9                    '%                     �    :                    H%                     �    ;                    i%                     �    <                    �%                     �    =                    �%                     5�_�  y  {          z  :       ����                                                                                                                                                                                                                                                                                                                M          1   9      5   :          :    f=     �  9  @  k           haso3 <= haso(127 downto 9);        haso4 <= haso(159 downto 1);        haso5 <= haso(191 downto 1);        haso6 <= haso(223 downto 1);        haso7 <= haso(255 downto 2);    �  :  ;  k    5��    9                    3%                     �    :                    V%                     �    ;                    y%                     �    <                    �%                     �    =                    �%                     5�_�  z  |          {  :       ����                                                                                                                                                                                                                                                                                                                M          1   9      5   :          :    f=     �  9  ;  k      "    haso3 <= haso(127 downto 96));5��    9                    4%                     5�_�  {  }          |  7       ����                                                                                                                                                                                                                                                                                                                M          1   9      5   :          :    f=   � �  6  8  k           haso0 <= haso(31 downto 0));5��    6                    �$                     5�_�  |  ~          }  .   ,    ����                                                                                                                                                                                                                                                                                                                M          1   9      5   :          :    f=.     �  -  /  k      ;    get_aout: adder32 port map (h0, av, haso(31 downto 0));5��    -  ,                  �"                     5�_�  }  �          ~  .   ,    ����                                                                                                                                                                                                                                                                                                                M          1   9      5   :          :    f=0     �  -  /  k      .    get_aout: adder32 port map (h0, av, haso);5��    -  ,                  �"                     5�_�  ~  �        �  /   ,    ����                                                                                                                                                                                                                                                                                                                M          1   9      5   :          :    f=:     �  3  5  k      >    get_gout: adder32 port map (h6, gv, haso(223 downto 192));�  2  4  k      >    get_fout: adder32 port map (h5, fv, haso(191 downto 160));�  1  3  k      >    get_eout: adder32 port map (h4, ev, haso(159 downto 128));�  0  2  k      =    get_dout: adder32 port map (h3, dv, haso(127 downto 96));�  /  1  k      <    get_cout: adder32 port map (h2, cv, haso(95 downto 64));�  .  0  k      <    get_bout: adder32 port map (h1, bv, haso(63 downto 32));5��    .  ,                 #                    �    /  ,                 M#                    �    0  ,                 }#                    �    1  ,                 �#                    �    2  ,                 �#                    �    3  ,                 $                    5�_�  �  �          �  5   ,    ����                                                                                                                                                                                                                                                                                                                M          1   9      5   :          :    f=<     �  4  6  k      >    get_hout: adder32 port map (hv, hv, haso(255 downto 224));5��    4  ,                  =$                     5�_�  �  �          �  5   ,    ����                                                                                                                                                                                                                                                                                                                M          1   9      5   :          :    f=>     �  4  6  k      .    get_hout: adder32 port map (hv, hv, haso);5��    4  ,                  =$                     5�_�  �  �          �  /   ,    ����                                                                                                                                                                                                                                                                                                                M          5   ,      /   ,          ,    f=B   � �  .  6  k      /    get_bout: adder32 port map (h1, bv, haso0);   /    get_cout: adder32 port map (h2, cv, haso0);   /    get_dout: adder32 port map (h3, dv, haso0);   /    get_eout: adder32 port map (h4, ev, haso0);   /    get_fout: adder32 port map (h5, fv, haso0);   /    get_gout: adder32 port map (h6, gv, haso0);   /    get_hout: adder32 port map (hv, hv, haso0);5��    .  ,                 #                    �    /  ,                 M#                    �    0  ,                 }#                    �    1  ,                 �#                    �    2  ,                 �#                    �    3  ,                 $                    �    4  ,                 =$                    5�_�  �  �          �  7       ����                                                                                                                                                                                                                                                                                                                M          7   
      7   
          
    f=\     �  6  8  k          haso0 <= haso(31 downto 0);5��    6                    F$                     5�_�  �  �          �  7       ����                                                                                                                                                                                                                                                                                                                M          7   
      7   
          
    f=b     �  6  8  k          <= haso(31 downto 0);5��    6                    Z$                     5�_�  �  �          �  7       ����                                                                                                                                                                                                                                                                                                                M          7   
      7   
          
    f=c     �  6  8  k          <= haso(31 downto 0) ;�  7  8  k    5��    6                    [$                     5�_�  �  �          �  7       ����                                                                                                                                                                                                                                                                                                                M          7   
      7   
          
    f=e     �  6  8  k           <= haso(31 downto 0) haso0 ;5��    6                    [$                     5�_�  �  �          �  7   "    ����                                                                                                                                                                                                                                                                                                                M          7   
      7   
          
    f=j     �  6  8  k      #    <= haso(31 downto 0) <= haso0 ;5��    6  !                  c$                     5�_�  �  �          �  7       ����                                                                                                                                                                                                                                                                                                                M          7   
      7   
          
    f=o     �  6  8  k      "    <= haso(31 downto 0) <= haso0;5��    6                    F$                     5�_�  �  �          �  8       ����                                                                                                                                                                                                                                                                                                                M          7   
      7   
          
    f=t     �  7  9  k           haso1 <= haso(63 downto 32);�  8  9  k    5��    7                    f$                     �    7                 
   {$              
       �    7  "                  �$                     �    7                    f$                     5�_�  �  �          �  9       ����                                                                                                                                                                                                                                                                                                                M          7   
      7   
          
    f=~   � �  =  ?  k      "    haso7 <= haso(255 downto 224);�  >  ?  k    �  <  >  k      "    haso6 <= haso(223 downto 192);�  =  >  k    �  ;  =  k      "    haso5 <= haso(191 downto 160);�  <  =  k    �  :  <  k      "    haso4 <= haso(159 downto 128);�  ;  <  k    �  9  ;  k      !    haso3 <= haso(127 downto 96);�  :  ;  k    �  8  :  k           haso2 <= haso(95 downto 64);�  9  :  k    5��    8                    �$                     �    8                 
   �$              
       �    8  "                  �$                     �    8                    �$                     �    9                    �$                     �    9                 
   �$              
       �    9  #                  �$                     �    9                    �$                     �    :                    �$                     �    :                 
   �$              
       �    :  $                  �$                     �    :                    �$                     �    ;                    �$                     �    ;                 
   %              
       �    ;  $                  %                     �    ;                    �$                     �    <                    %                     �    <                 
   '%              
       �    <  $                  0%                     �    <                    %                     �    =                    3%                     �    =                 
   J%              
       �    =  $                  S%                     �    =                    3%                     5�_�  �  �          �  U       ����                                                                                                                                                                                                                                                                                                                M                                            fB�
     �  T  V  k      '    current_w <= w_vec(511 downto 480);5��    T                   �&                    �    T                    �&                     5�_�  �  �          �  U   !    ����                                                                                                                                                                                                                                                                                                                M                                            fB�   � �  T  V  k      &    current_w <= w_vec(31 downto 480);5��    T  !                 �&                    5�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                M                                            fB��     �   3   5  k      2            vector <= vector(479 downto 0) & data;5��    3                    T                    5�_�  �  �          �   4   -    ����                                                                                                                                                                                                                                                                                                                M                                            fB��     �   3   5  k      2            vector <= vector(511 downto 0) & data;5��    3   -                  d                     5�_�  �  �  �      �   4       ����                                                                                                                                                                                                                                                                                                                M                                            fB��     �   3   5  k      .            vector <= vector(511 downto 0) & ;�   4   5  k    5��    3                     M                     5�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                M                                            fB��     �   3   5  k      2            vector <= datavector(511 downto 0) & ;5��    3                     Q                     5�_�  �  �          �   4   1    ����                                                                                                                                                                                                                                                                                                                M                                            fB��     �   3   5  k      5            vector <= data & vector(511 downto 0) & ;5��    3   1                  h                     5�_�  �  �          �   4   1    ����                                                                                                                                                                                                                                                                                                                M                                            fB��     �   3   5  k      4            vector <= data & vector(511 downto 0)& ;5��    3   1                  h                     5�_�  �  �          �   4   /    ����                                                                                                                                                                                                                                                                                                                M                                            fB��   � �   3   5  k      2            vector <= data & vector(511 downto 0);5��    3   /                 f                    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                M                                            fB��     �      k      <    int1: sigma1 port map(w_vec(63 downto 32), op1); -- t-145��                        �                    5�_�  �  �          �     +    ����                                                                                                                                                                                                                                                                                                                M                                            fB��     �      k      =    int1: sigma1 port map(w_vec(479 downto 32), op1); -- t-145��      +                 �                    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                M                                            fB�     �      k      =    int2: sigma0 port map(w_vec(479 downto 448), op2); -- t-15��                        �                    5�_�  �  �          �     *    ����                                                                                                                                                                                                                                                                                                                M                                            fB�     �      k      <    int2: sigma0 port map(w_vec(63 downto 448), op2); -- t-15��      *                 �                    5�_�  �  �          �     <    ����                                                                                                                                                                                                                                                                                                                M                                            fB�L     �      k      >    int1: sigma1 port map(w_vec(479 downto 448), op1); -- t-145��      <                 �                    5�_�  �  �          �     :    ����                                                                                                                                                                                                                                                                                                                M                                            fB�Q     �      k      ;    int2: sigma0 port map(w_vec(63 downto 32), op2); -- t-15��      :                 �                    5�_�  �  �          �     T    ����                                                                                                                                                                                                                                                                                                                M                                            fB�Z     �      k      [    int3: adder32 port map(w_vec(223 downto 192), w_vec(511 downto 480), op4); -- t-9 and t5��      T                 z                    5�_�  �  �          �     [    ����                                                                                                                                                                                                                                                                                                                M                                            fB�`     �      k      [    int3: adder32 port map(w_vec(223 downto 192), w_vec(511 downto 480), op4); -- t-7 and t5��      [                  �                     5�_�  �  �          �     !    ����                                                                                                                                                                                                                                                                                                                M                                            fB�i     �      k      ^    int3: adder32 port map(w_vec(223 downto 192), w_vec(511 downto 480), op4); -- t-7 and t-165��      !                 G                    5�_�  �  �          �     ,    ����                                                                                                                                                                                                                                                                                                                M                                            fB�o     �      k      ^    int3: adder32 port map(w_vec(319 downto 192), w_vec(511 downto 480), op4); -- t-7 and t-165��      ,                 R                    5�_�  �  �          �     8    ����                                                                                                                                                                                                                                                                                                                M                                            fB�y     �      k      ^    int3: adder32 port map(w_vec(319 downto 288), w_vec(511 downto 480), op4); -- t-7 and t-165��      8                 ^                    5�_�  �  �          �     B    ����                                                                                                                                                                                                                                                                                                                M                                            fB�{   � �      k      ]    int3: adder32 port map(w_vec(319 downto 288), w_vec(31 downto 480), op4); -- t-7 and t-165��      B                 h                    �      B                 h                    5�_�  �              �  5   !    ����                                                                                                                                                                                                                                                                                                                M                                            fB�   � �  4  6  k      /    get_hout: adder32 port map (hv, hv, haso7);5��    4  !                 3$                    5�_�  �          �  �   4       ����                                                                                                                                                                                                                                                                                                                M                                            fB��     �   4   5  k    �   3   5  k      2            vector <= vdataector(511 downto 0) & ;5��    3                     N                     5�_�  ~          �    /   ,    ����                                                                                                                                                                                                                                                                                                                M          1   9      5   :          :    f=6     �  .  0  k      /    get_bout: adder32 port map (h1, bv, haso0);�  /  1  k      /    get_cout: adder32 port map (h2, cv, haso0);�  0  2  k      /    get_dout: adder32 port map (h3, dv, haso0);�  1  3  k      /    get_eout: adder32 port map (h4, ev, haso0);�  2  4  k      /    get_fout: adder32 port map (h5, fv, haso0);�  3  5  k      /    get_gout: adder32 port map (h6, gv, haso0);�  4  6  k      !    get_hout: adder32 port map 0;5��    .  ,                 #                    �    /  ,                 M#                    �    0  ,                 }#                    �    1  ,                 �#                    �    2  ,                 �#                    �    3  ,                 $                    �    4                   0$                    5�_�  v          x  w  8       ����                                                                                                                                                                                                                                                                                                                M          8         >                 f=�     �  7  ?  k          haso-1 <= haso();       haso-1 <= haso();       haso-1 <= haso();       haso-1 <= haso();       haso-1 <= haso();       haso-1 <= haso();       haso-1 <= haso();5��    7                   �$                    �    8                   �$                    �    9                   �$                    �    :                   %                    �    ;                   '%                    �    <                   =%                    �    =                   S%                    5�_�  o          q  p  6        ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=�     �  6  7  c    �  5  ?  c   	   haso0   haso1   !haso2    step: stepfun port map (   haso3        ai => a_reg,   haso4        bi => b_reg,   haso5        ci => c_reg,   haso6        di => d_reg,   haso7        ei => e_reg,           fi => f_reg,5��    5                     �$                     �    6                     �$                     �    7                     �$                     �    8                     �$                     �    9                     �$                     �    :                     %                     �    ;                     -%                     �    <                     G%                     5�_�  d      f  h  g   �       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=%     �   �   �  b      *    signal haso1: bit_vector(31 downto 0);   *    signal haso1: bit_vector(31 downto 0);   *    signal haso1: bit_vector(31 downto 0);   *    signal haso1: bit_vector(31 downto 0);   *    signal haso1: bit_vector(31 downto 0);   *    signal haso1: bit_vector(31 downto 0);   *    signal haso1: bit_vector(31 downto 0);5��    �                    V                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                                        �    �                    -                    �    �                    X                    5�_�  d      e  g  f   �       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=!     �   �   �  b      )    signal haso: bit_vector(31 downto 0);   *    signal hasoa: bit_vector(31 downto 0);   *    signal hasoa: bit_vector(31 downto 0);   *    signal hasoa: bit_vector(31 downto 0);   *    signal hasoa: bit_vector(31 downto 0);   *    signal hasoa: bit_vector(31 downto 0);   *    signal hasoa: bit_vector(31 downto 0);�   �   �  b      *    signal hasoa: bit_vector(31 downto 0);5��    �                     V                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     (                     �    �                     R                     �    �                     V                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                                          �    �                     -                     �    �                     X                     5�_�  d          f  e   �       ����                                                                                                                                                                                                                                                                                                                M           �          �                 f=     �   �   �  b      *    signal haso1: bit_vector(31 downto 0);   *    signal haso1: bit_vector(31 downto 0);   *    signal haso1: bit_vector(31 downto 0);   *    signal haso1: bit_vector(31 downto 0);   *    signal haso1: bit_vector(31 downto 0);   *    signal haso1: bit_vector(31 downto 0);   *    signal haso1: bit_vector(31 downto 0);5��    �                    V                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                                        �    �                    -                    �    �                    X                    5�_�  ^  `      d  _   �   )    ����                                                                                                                                                                                                                                                                                                                M                                            f=
     �   �   �  [    �   �   �  [      *    signal haso0: bit_vector(31 downto 0);5��    �                      G              +       5�_�  _  a          `   �       ����                                                                                                                                                                                                                                                                                                                M                                            f=     �   �   �  \    �   �   �  \      *    signal haso0: bit_vector(31 downto 0);5��    �                      r              +       5�_�  `  b          a   �       ����                                                                                                                                                                                                                                                                                                                M                                            f=     �   �   �  ]    �   �   �  ]      *    signal haso0: bit_vector(31 downto 0);5��    �                      �              +       5�_�  a  c          b   �       ����                                                                                                                                                                                                                                                                                                                M                                            f=     �   �   �  ^    �   �   �  ^      *    signal haso0: bit_vector(31 downto 0);5��    �                      �              +       5�_�  b              c   �       ����                                                                                                                                                                                                                                                                                                                M                                            f=     �   �   �  _    �   �   �  _      *    signal haso0: bit_vector(31 downto 0);5��    �                      �              +       5�_�  
             <        ����                                                                                                                                                                                                                                                                                                                N           <          <          V       f(A/     �   ;   [        5��    ;                      �      �              5�_�                 <        ����                                                                                                                                                                                                                                                                                                                M           <          <          V       f(A0   � �   ;   =        5��    ;                      �                     5�_�                 d       ����                                                                                                                                                                                                                                                                                                                M           <          <          V       f(AZ     �   c   e  9      !    component counter_generic  is5��    c                    �                    5�_�                 f       ����                                                                                                                                                                                                                                                                                                                M           <          <          V       f(Ag     �   e   g  9      N            clk, rst, start: in bit;                            -- Clock input5��    e                     �                     5�_�                 h       ����                                                                                                                                                                                                                                                                                                                M           i   	       e          V       f(Ar     �   g   i  9      F            count : out natural       -- 6-bit count output (64 steps)5��    g                    i	                    5�_�                 e       ����                                                                                                                                                                                                                                                                                                                M           e          l                 f(A}     �   d   j        �   e   f  4    �   d   e  4          generic(           MAX_COUNT: natural       );   
    port (   J        clk, rst, start: in bit;                            -- Clock input           done: out bit;   B        count : out natural       -- 6-bit count output (64 steps)       );5��    d                      �      �               �    d                      �              �       5�_�                 e       ����                                                                                                                                                                                                                                                                                                                M                                            f(A�   � �   d   f  <              generic(�   e   m  <                  MAX_COUNT: natural   
        );           port (   N            clk, rst, start: in bit;                            -- Clock input               done: out bit;   F            count : out natural       -- 6-bit count output (64 steps)   
        );5��    d                     �                     �    e                     �                     �    f                     	                     �    g                     	                     �    h                     &	                     �    i                     u	                     �    j                     �	                     �    k                     �	                     5�_�                 �       ����                                                                                                                                                                                                                                                                                                                M                                            f(A�     �   �   �  <      C    counter: counter_generic port map (clk, rst, ended, iteration);5��    �                    i                    �    �                     m                     �    �                     l                     �    �                     k                     �    �                     j                     �    �                 	   i             	       �    �                     q                     �    �                     p                     �    �                     o                     �    �                     n                     �    �                     m                     �    �                     l                     �    �                     k                     �    �                     j                     �    �                    i                    �    �                     w                     �    �                     v                     �    �                     u                     �    �                     t                     �    �                     s                     �    �                     r                     �    �                     q                     �    �                     p                     �    �                     o                     �    �                     n                     �    �                     m                     �    �                     l                     �    �                     k                     �    �                     j                     �    �                    i                    �    �                    i                    �    �                    i                    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                M                                            f(A�     �   �   �  <          counter: counter_generic    *    port map (clk, rst, ended, iteration);5��    �                    y                     5�_�                 �       ����                                                                                                                                                                                                                                                                                                                M                                            f(A�     �   �   �  =      .        port map (clk, rst, ended, iteration);5��    �                     ~                     5�_�                 �       ����                                                                                                                                                                                                                                                                                                                M                                            f(A�     �   �   �  =          �   �   �  >              generic map5��    �                      z              	       �    �                     z                    �    �                    �                    �    �                    �                    �    �                    �                    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                M                                            f(A�     �   �   �  >              generic map()5��    �                     �                     5�_�                 �       ����                                                                                                                                                                                                                                                                                                                M                                            f(A�     �   �   �  >              generic map(64)5��    �                     �                     5�_�                 �       ����                                                                                                                                                                                                                                                                                                                M                                            f(A�     �   �   �  >          signal iteration: natural;5��    �                    f                    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                M                                            f(A�     �   �   �  >          �   �   �  ?          signal enable;5��    �                      o                     �    �                     s                     5�_�                 �       ����                                                                                                                                                                                                                                                                                                                M                                            f(A�     �   �   �  ?          signal enable: bit;5��    �                     �                     5�_�                        ����                                                                                                                                                                                                                                                                                                                M                                            f(B     �   �    ?      6        port map (clk, rst, enable, ended, iteration);5��    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�              *       ����                                                                                                                                                                                                                                                                                                                M                                            f(Be     �  )  +  ?      &    current_k <= k_const((iteration));5��    )         
           �"      
               5�_�                 *       ����                                                                                                                                                                                                                                                                                                                M                                            f(Be     �  )  +  ?      %    current_k <= k_const(iteration));5��    )                    �"                     5�_�    !             *   "    ����                                                                                                                                                                                                                                                                                                                M                                            f(Bf   � �  )  +  ?      $    current_k <= k_const(iteration);5��    )  "                  �"                     5�_�     "          !  &        ����                                                                                                                                                                                                                                                                                                                M           e          l                 f(B�     �  &  '  ?       5��    &                     f"                     �    &                     f"                     5�_�  !  #          "  '        ����                                                                                                                                                                                                                                                                                                                M           e          l                 f(B�     �  '  (  @    �  '  (  @          process(clk, rst)   	    begin           if rst = '0' then               enable <= '1';           end if;           if rst = '1' then               done <= '0';               enable <= '0';   #        elsif rising_edge(clk) then   "            if iteration = 63 then                   done <= '1';               end if;               -- Update kpw   (        current_k <= k_const(iteration);   +        current_w <= w_vec(511 downto 480);           end if;               end process;5��    '                     g"              �      5�_�  "  $          #  :        ����                                                                                                                                                                                                                                                                                                                M          7         5          V       f(B�     �  9  ;        5��    9                     $                     5�_�  #  %          $  5       ����                                                                                                                                                                                                                                                                                                                M          (         7          V       f(B�     �  4  8        5��    4                     �#      k               5�_�  $  )          %  7       ����                                                                                                                                                                                                                                                                                                                M          (         7          V       f(B�     �  '  8  P          -- process(clk, rst)       -- begin       --     if rst = '0' then       --         enable <= '1';       --     end if;       --     if rst = '1' then       --         done <= '0';       --         enable <= '0';   &    --     elsif rising_edge(clk) then   %    --         if iteration = 63 then       --             done <= '1';       --         end if;       --       --     end if;       --       -- end process;5��    '                    g"      N      �      5�_�  %  *  &      )  7       ����                                                                                                                                                                                                                                                                                                                M          (         7          V       f(Cz     �  '  8  P          process(clk, rst)   	    begin           if rst = '0' then               enable <= '1';           end if;           if rst = '1' then               done <= '0';               enable <= '0';   #        elsif rising_edge(clk) then   "            if iteration = 63 then                   done <= '1';               end if;               end if;           end process;5��    '                    g"      �      N      5�_�  )  +          *  2       ����                                                                                                                                                                                                                                                                                                                M          (         7          V       f(C�     �  1  3  P                      enable <= '1';5��    1                   q#                    5�_�  *  ,          +  2       ����                                                                                                                                                                                                                                                                                                                M          *         ,          V       f(C�     �  1  3  P                      enable <= '0';5��    1                   |#                    5�_�  +  -          ,  *        ����                                                                                                                                                                                                                                                                                                                M          *         *          V       f(C�     �  )  -        5��    )                     �"      E               5�_�  ,  .          -  +       ����                                                                                                                                                                                                                                                                                                                M          *         *          V       f(C�     �  *  ,        5��    *                     �"                     5�_�  -  /          .  +       ����                                                                                                                                                                                                                                                                                                                M          *         *          V       f(C�     �  *  ,  L                  enable <= '1';5��    *                   �"                    5�_�  .  0          /  +       ����                                                                                                                                                                                                                                                                                                                M          *         *          V       f(C�     �  *  ,  L                  enable <= '0';5��    *                   �"                    5�_�  /  1          0  +       ����                                                                                                                                                                                                                                                                                                                M          *         *          V       f(C�     �  *  ,  L                  enable <= '1';5��    *                   �"                    5�_�  0  2          1   A       ����                                                                                                                                                                                                                                                                                                                M          *         *          V       f(D>     �   @   B  L      "        clk, rst, enable : in bit;5��    @                                          5�_�  1  3          2   A       ����                                                                                                                                                                                                                                                                                                                M          *         *          V       f(DB     �   @   B  L      !        clk, rst, enable: in bit;5��    @                                          5�_�  2  4          3   �       ����                                                                                                                                                                                                                                                                                                                M          '         2          V       f(DK     �   �   �        5��    �                      v                     5�_�  3  5          4  2       ����                                                                                                                                                                                                                                                                                                                M          
   %         %          %    f(D�   � �  &  3  K          -- process(clk, rst)       -- begin       --     if rst = '1' then       --         enable <= '1';   &    --     elsif rising_edge(clk) then   %    --         if iteration = 63 then   !    --             enable <= '0';       --         end if;       --       --     end if;       --       -- end process;5��    &                    V"      �             5�_�  4  6          5  
   &    ����                                                                                                                                                                                                                                                                                                                M             %         %          %    f(G>     �  	    K      >    get_aout: adder32 port map (h0, a_reg, haso(31 downto 0));�  
    K      ?    get_bout: adder32 port map (h1, bvreg, haso(63 downto 32));   ?    get_cout: adder32 port map (h2, cvreg, haso(95 downto 64));   @    get_dout: adder32 port map (h3, dvreg, haso(127 downto 96));   A    get_eout: adder32 port map (h4, evreg, haso(159 downto 128));   A    get_fout: adder32 port map (h5, fvreg, haso(191 downto 160));   A    get_gout: adder32 port map (h6, gvreg, haso(223 downto 192));   A    get_hout: adder32 port map (hv, hvreg, haso(255 downto 224));5��    	  %                                     �    
  &                  R                     �      &                  �                     �      &                  �                     �      &                                        �      &                  U                      �      &                  �                      �      &                  �                      5�_�  5  7          6     %    ����                                                                                                                                                                                                                                                                                                                M          
   %         (          (    f(GC   � �  
    K      ?    get_bout: adder32 port map (h1, b_reg, haso(63 downto 32));   ?    get_cout: adder32 port map (h2, c_reg, haso(95 downto 64));   @    get_dout: adder32 port map (h3, d_reg, haso(127 downto 96));   A    get_eout: adder32 port map (h4, e_reg, haso(159 downto 128));   A    get_fout: adder32 port map (h5, f_reg, haso(191 downto 160));   A    get_gout: adder32 port map (h6, g_reg, haso(223 downto 192));   A    get_hout: adder32 port map (hv, h_reg, haso(255 downto 224));5��    
  %                 Q                    �      %                 �                    �      %                 �                    �      %                                      �      %                 T                     �      %                 �                     �      %                 �                     5�_�  6  9          7  
   %    ����                                                                                                                                                                                                                                                                                                                M          
   %         %          %    f(H   � �  	    K      :    get_aout: adder32 port map (h0, a, haso(31 downto 0));   <    get_bout: adder32 port map (h1, bv, haso(63 downto 32));   <    get_cout: adder32 port map (h2, cv, haso(95 downto 64));   =    get_dout: adder32 port map (h3, dv, haso(127 downto 96));   >    get_eout: adder32 port map (h4, ev, haso(159 downto 128));   >    get_fout: adder32 port map (h5, fv, haso(191 downto 160));   >    get_gout: adder32 port map (h6, gv, haso(223 downto 192));   >    get_hout: adder32 port map (hv, hv, haso(255 downto 224));�  	    K      ;    get_aout: adder32 port map (h0, av, haso(31 downto 0));5��    	  %                                       �    
  %                  M                     �      %                  �                     �      %                  �                     �      %                                        �      %                  @                      �      %                  ~                      �      %                  �                      �    	  %                                       �    
  %                  N                     �      %                  �                     �      %                  �                     �      %                                        �      %                  E                      �      %                  �                      �      %                  �                      5�_�  7  :  8      9  
   &    ����                                                                                                                                                                                                                                                                                                                M             %         %          %    f(I�     �  	    K      >    get_aout: adder32 port map (h0, a_reg, haso(31 downto 0));�  
    K      ?    get_bout: adder32 port map (h1, bvreg, haso(63 downto 32));   ?    get_cout: adder32 port map (h2, cvreg, haso(95 downto 64));   @    get_dout: adder32 port map (h3, dvreg, haso(127 downto 96));   A    get_eout: adder32 port map (h4, evreg, haso(159 downto 128));   A    get_fout: adder32 port map (h5, fvreg, haso(191 downto 160));   A    get_gout: adder32 port map (h6, gvreg, haso(223 downto 192));   A    get_hout: adder32 port map (hv, hvreg, haso(255 downto 224));5��    	  %                                     �    
  &                  R                     �      &                  �                     �      &                  �                     �      &                                        �      &                  U                      �      &                  �                      �      &                  �                      5�_�  9  ;          :     %    ����                                                                                                                                                                                                                                                                                                                M          '         2          V   %    f(I�   � �  
    K      ?    get_bout: adder32 port map (h1, b_reg, haso(63 downto 32));   ?    get_cout: adder32 port map (h2, c_reg, haso(95 downto 64));   @    get_dout: adder32 port map (h3, d_reg, haso(127 downto 96));   A    get_eout: adder32 port map (h4, e_reg, haso(159 downto 128));   A    get_fout: adder32 port map (h5, f_reg, haso(191 downto 160));   A    get_gout: adder32 port map (h6, g_reg, haso(223 downto 192));   A    get_hout: adder32 port map (hv, h_reg, haso(255 downto 224));5��    
  %                 Q                    �      %                 �                    �      %                 �                    �      %                                      �      %                 T                     �      %                 �                     �      %                 �                     5�_�  :  <          ;  2       ����                                                                                                                                                                                                                                                                                                                M          '         2          V   %    f(N�     �  &  3  K          process(clk, rst)   	    begin           if rst = '1' then               enable <= '1';   #        elsif rising_edge(clk) then   "            if iteration = 63 then                   enable <= '0';               end if;               end if;           end process;5��    &                    n"            �       5�_�  ;  =          <  +       ����                                                                                                                                                                                                                                                                                                                M          '         2          V   %    f(N�     �  *  ,  K      $            if rising_edge(clk) then5��    *                   �"                    �    *                    �"                    5�_�  <  >          =  ,       ����                                                                                                                                                                                                                                                                                                                M          '         2          V   %    f(N�     �  +  -  K      &                if iteration = 63 then5��    +                    �"                     5�_�  =  ?          >  4       ����                                                                                                                                                                                                                                                                                                                M          '         2          V   %    f(N�     �  3  5        5��    3                     f#                     5�_�  >  @          ?  -       ����                                                                                                                                                                                                                                                                                                                M          '         2          V   %    f(N�     �  ,  .  J                      done <= '0';5��    ,                   #                    5�_�  ?  A          @  *       ����                                                                                                                                                                                                                                                                                                                M          '         2          V   %    f(N�     �  )  +  J                  done <= '1';5��    )                   �"                    5�_�  @  B          A  -       ����                                                                                                                                                                                                                                                                                                                M          '         2          V   %    f(N�     �  ,  .  J                           done <= '0';5��    ,                    #                     5�_�  A  G          B  -       ����                                                                                                                                                                                                                                                                                                                M          '         3          V   %    f(N�   � �  -  .  J                          �  -  /  K                      end if;5��    -                     .#                     �    -                    B#                     �    -                    .#                    �    -                    B#                     5�_�  B  H  C      G  '       ����                                                                                                                                                                                                                                                                                                                M          '         3          V   %    f(O@   � �  &  (  K          process(clk, rst, enable)5��    &                    �"                     �    &                    �"                     �    &                    �"                     �    &                   �"                    �    &                   �"                    �    &                    �"                     �    &                   �"                    5�_�  G  I          H  ,        ����                                                                                                                                                                                                                                                                                                                M          '         3          V   %    f(OX   � �  +  -  K      &                if iteration = 62 then5��    +                    #                    5�_�  H  J          I  +       ����                                                                                                                                                                                                                                                                                                                M          '         3          V   %    f(Ol     �  *  ,  K      '            elsif rising_edge(clk) then5��    *                    �"                     5�_�  I  K          J  +       ����                                                                                                                                                                                                                                                                                                                M          '         3          V   %    f(Oo     �  *  ,  K      #        elsif rising_edge(clk) then5��    *                    �"                     5�_�  J  L          K  ,       ����                                                                                                                                                                                                                                                                                                                M          ,         ,          v       f(Ot     �  +  -  K      #                iteration = 62 then5��    +                    �"                     5�_�  K  M          L  ,       ����                                                                                                                                                                                                                                                                                                                M          ,         ,          v       f(Oz     �  +  -  K                       then5��    +                    �"                     5�_�  L  N          M  +       ����                                                                                                                                                                                                                                                                                                                M          ,         ,          v       f(O|     �  *  ,  K      $        elsif rising_edge(clk)  then5��    *                    �"                     5�_�  M  O          N  +       ����                                                                                                                                                                                                                                                                                                                M          ,         ,          v       f(O}     �  +  ,  K    �  *  ,  K      2        elsif rising_edge(clk) iteration = 62 then5��    *                    �"                     5�_�  N  P          O  +   ,    ����                                                                                                                                                                                                                                                                                                                M          ,         ,          v       f(O     �  *  ,  K      2        elsif rising_edge(clk) iteration = 63 then5��    *  ,                 �"                    5�_�  O  Q          P  +       ����                                                                                                                                                                                                                                                                                                                M          ,         ,          v       f(O�     �  *  ,  K      6        elsif rising_edge(clk) and iteration = 63 then5��    *                    �"                     5�_�  P  R          Q  ,       ����                                                                                                                                                                                                                                                                                                                M          ,         ,          v       f(O�     �  +  -        5��    +                      #                     5�_�  Q  S          R  -       ����                                                                                                                                                                                                                                                                                                                M          ,         ,          v       f(O�     �  ,  .        5��    ,                     !#                     5�_�  R  T          S  ,       ����                                                                                                                                                                                                                                                                                                                M          ,         ,          v       f(O�     �  +  -  I                      done <= '0';5��    +                    #                     5�_�  S  U          T  -       ����                                                                                                                                                                                                                                                                                                                M          ,         ,          v       f(O�     �  ,  .  I              end if;5��    ,                    %#                     5�_�  T  V          U  /       ����                                                                                                                                                                                                                                                                                                                M          ,         ,          v       f(O�     �  .  0        5��    .                     .#                     5�_�  U  W          V  .        ����                                                                                                                                                                                                                                                                                                                M          ,         ,          v       f(O�   � �  -  /        5��    -                     -#                     5�_�  V  X          W  ,       ����                                                                                                                                                                                                                                                                                                                M          '         /          V       f(O�     �  +  -  G                  done <= '0';5��    +                    #                     5�_�  W  Y          X  /       ����                                                                                                                                                                                                                                                                                                                M          '         /          V       f(g�     �  &  0  G   	        -- process(clk, rst, enable)       -- begin       --     if rst = '1' then       --         done <= '1';   9    --     elsif rising_edge(clk) and iteration = 63 then       --         done <= '0';       --     end if;       --       -- end process;5��    &      	       	       n"      �       �       5�_�  X              Y  0        ����                                                                                                                                                                                                                                                                                                                M          '         /          V       f(g�     �  0  1  G          �  0  2  H          done <= ended;5��    0                     Z#                     �    0                     Z#                     �    0                    e#                     �    0  
                 d#                    �    0                    i#                     �    0                    h#                     �    0                    g#                     �    0                   f#                    �    0                   f#                    �    0                   f#                    5�_�  B  D      G  C  +       ����                                                                                                                                                                                                                                                                                                                M          '         3          V   %    f(O     �  *  ,  K      7            if rising_edge(clk) and iteration = 63 then5��    *                    �"                     �    *  &                  �"                     �    *  %                  �"                     �    *  $              	   �"             	       �    *  $       	          �"      	              �    *  $                 �"                    5�_�  C  E          D  ,   %    ����                                                                                                                                                                                                                                                                                                                M          '         2          V   %    f(O     �  +  -        5��    +                     �"      '               5�_�  D  F          E  ,       ����                                                                                                                                                                                                                                                                                                                M          '         2          V   %    f(O     �  +  -  J                      done <= '0';5��    +                    #                     �    +                    	#                     5�_�  E              F  -       ����                                                                                                                                                                                                                                                                                                                M          '         1          V   %    f(O   � �  ,  .        5��    ,                     #                     5�_�  7          9  8   �       ����                                                                                                                                                                                                                                                                                                                M          
   %         (          (    f(H�   � �   �   �  K              generic map(63)5��    �                    �                    5�_�  %  '      )  &          ����                                                                                                                                                                                                                                                                                                                M          (         7          V       f(B�     �   �    P      0        port map (clk, rst, , ended, iteration);5��    �                     �                     5�_�  &  (          '          ����                                                                                                                                                                                                                                                                                                                M          (         7          V       f(B�     �   �    P      2        port map (clk, rst, '', ended, iteration);5��    �                     �                     5�_�  '              (          ����                                                                                                                                                                                                                                                                                                                M          (         7          V       f(B�   � �   �    P      3        port map (clk, rst, '1', ended, iteration);5��    �                     �                     5�_�                *       ����                                                                                                                                                                                                                                                                                                                M                                            f(Bb     �  )  +  ?      )    current_k <= (to_integer(iteration));5��    )                    �"                     5�_�  �           �   V       ����                                                                                                                                                                                                                                                                                                                l           V   
       V          V       f�     �   U   Y        5��    U                             T               5�_�  �                  I        ����                                                                                                                                                                                                                                                                                                                o           Y   
       Y          V       f�     �   I   J  X    �   I   J  X      2    if rst = '0' and to_integer(counter) = 63 then           done <= '1';       end if;5��    I                                    T       5�_�  �          �  �   W       ����                                                                                                                                                                                                                                                                                                                m           W          V          V       f     �   V   Y        �   U   W  Y       5��    V                      c      2               �    U          >           $      >               �    U                     #                     �    U                     "                     �    U                     !                     �    U                                            5�_�  �  �      �  �   R        ����                                                                                                                                                                                                                                                                                                                l           R   (       R          V   (    f)     �   Q   U        5��    Q                      �      [               5�_�  �  �          �   U       ����                                                                                                                                                                                                                                                                                                                m           R   (       R          V   (    f.     �   U   V  X       5��    U                      7                     �    U                      7                     5�_�  �  �          �   V        ����                                                                                                                                                                                                                                                                                                                p           W          Y                 f/     �   V   W  Y    �   V   W  Y      ,            if to_integer(counter) = 63 then                   done <= '1';               else5��    V                      8              [       5�_�  �  �          �   W       ����                                                                                                                                                                                                                                                                                                                p           W          Y                 f2     �   V   X  \      $    if to_integer(counter) = 63 then5��    V                     <                     5�_�  �  �          �   X       ����                                                                                                                                                                                                                                                                                                                p           W          Y                 f3     �   W   Y  \              done <= '1';5��    W                    a                    5�_�  �  �          �   Y       ����                                                                                                                                                                                                                                                                                                                p           W          Y                 f5     �   X   Z  \          else5��    X                     v                     5�_�  �  �          �   Y       ����                                                                                                                                                                                                                                                                                                                p           W          Y                 f7     �   X   Z  \          end if.5��    X                    v                    5�_�  �  �          �   Y   
    ����                                                                                                                                                                                                                                                                                                                p           W          Y                 f:     �   X   Z  \          end if;5��    X   
                 |                    5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                p           W          Y                 fB     �   R   T  \              end if;5��    R                                          5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                o           V          X                 fC     �   R   T        5��    R                      �                     5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                o           V          X                 fE     �   Q   S  [      #            counter <= counter + 1;5��    Q                     �                     5�_�  �  �          �   V       ����                                                                                                                                                                                                                                                                                                                o           V          X                 fd     �   U   W  [      -    generate if to_integer(counter) = 63 then5��    U                  	   $              	       5�_�  �              �   V       ����                                                                                                                                                                                                                                                                                                                o                                            fi   � �   U   W  [      $    if to_integer(counter) = 63 then5��    U          	           $      	               5�_�  �          �  �  '   %    ����                                                                                                                                                                                                                                                                                                                o          '   %      .   %          %    f=   � �  &  /  [      :    get_aout: adder32 port map (h0, a, haso(31 downto 0));   ?    get_bout: adder32 port map (h1, b_reg, haso(63 downto 32));   ?    get_cout: adder32 port map (h2, c_reg, haso(95 downto 64));   @    get_dout: adder32 port map (h3, d_reg, haso(127 downto 96));   A    get_eout: adder32 port map (h4, e_reg, haso(159 downto 128));   A    get_fout: adder32 port map (h5, f_reg, haso(191 downto 160));   A    get_gout: adder32 port map (h6, g_reg, haso(223 downto 192));   A    get_hout: adder32 port map (hv, h_reg, haso(255 downto 224));�  &  (  [      >    get_aout: adder32 port map (h0, a_reg, haso(31 downto 0));5��    &  %                  �!                     �    '  %                  �!                     �    (  %                  2"                     �    )  %                  n"                     �    *  %                  �"                     �    +  %                  �"                     �    ,  %                  '#                     �    -  %                  e#                     �    &  %                  �!                     �    '  %                  �!                     �    (  %                  :"                     �    )  %                  z"                     �    *  %                  �"                     �    +  %                  �"                     �    ,  %                  ?#                     �    -  %                  �#                     5�_�  �          �  �   �       ����                                                                                                                                                                                                                                                                                                                o           �          �          v       f     �   �   �  m          signal ended: bit;5��    �                     M                     5�_�  �          �  �   R       ����                                                                                                                                                                                                                                                                                                                o          &   %      -   (          (    f �     �   Q   S  m      -            if counter = to_unsigned(63) then5��    Q                     �                     5�_�  �  �      �  �          ����                                                                                                                                                                                                                                                                                                                i              %      '   (          (    f      �        g               rst, clk enable: in bit;5��                         T                      5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                i              %      '   (          (    f      �        g              rst, clkenable: in bit;5��                         T                      5�_�  �              �          ����                                                                                                                                                                                                                                                                                                                i              %      '   (          (    f      �        g              rst, clk: in bit;5��                         T                      5�_�  �  �      �  �  >       ����                                                                                                                                                                                                                                                                                                                i          !   %      (   (          (    f�f     �  =  ?  h          process(, rst)5��    =                    �$                     5�_�  �  �          �  >       ����                                                                                                                                                                                                                                                                                                                i          !   %      (   (          (    f�g     �  =  ?  h          process(rst)5��    =                    �$                     5�_�  �  �          �  C       ����                                                                                                                                                                                                                                                                                                                i          !   %      (   (          (    f�o     �  B  D  h              els then5��    B                    �$                     5�_�  �  �          �  C       ����                                                                                                                                                                                                                                                                                                                i          !   %      (   (          (    f�p     �  B  D  h              else then5��    B                    �$                     5�_�  �  �          �  C       ����                                                                                                                                                                                                                                                                                                                i          !   %      (   (          (    f�r     �  B  D  h              else 5��    B                    �$                     5�_�  �              �  C       ����                                                                                                                                                                                                                                                                                                                i          !   %      (   (          (    f�r   � �  B  D  h              else5��    B                    �$                     5�_�  �          �  �     6    ����                                                                                                                                                                                                                                                                                                                i           �          �   *       v   *    f��     �            5��                         �      B               5�_�  `  b      f  a     9    ����                                                                                                                                                                                                                                                                                                                i          P         T           V   9    f�     �      n      O    -- get_k: reg32 port map (rst, clk, enable, k_const(0), next_k, current_k);5��                        �      M       P       5�_�  a  c          b  Q        ����                                                                                                                                                                                                                                                                                                                i          P         Q           V   9    f�     �  P  U        �  O  Q  j                   current_k <= k_const5��    P                     �&      i               �    O                   x&                    �    O                    z&                     �    O                    y&                     �    O                	   x&             	       �    O         	          x&      	              �    O                   x&                    �    O                    �&                     �    O                    �&                     �    O                   �&                    �    O                   �&                    �    O                   �&                    5�_�  b  d          c  P        ����                                                                                                                                                                                                                                                                                                                i          P         Q           V   9    f�     �  O  Q  j      "            current_k <= k_const()5��    O                     �&                     5�_�  c  e          d  P   !    ����                                                                                                                                                                                                                                                                                                                i          P         Q           V   9    f�     �  O  Q  j      +            current_k <= k_const(iteration)5��    O  !                  �&                     �    O  !              	   �&             	       �    O  !       	          �&      	              �    O  !              	   �&             	       5�_�  d              e  P   +    ����                                                                                                                                                                                                                                                                                                                i          P         Q           V   9    f�   � �  O  Q  j      ,            current_k <= k_const(iteration);5��    O  +                  �&                     5�_�  0  2      =  1          ����                                                                                                                                                                                                                                                                                                                i          K         K   "       V   '    f�   � �            5��                         �      N               5�_�  1  3          2  M       ����                                                                                                                                                                                                                                                                                                                i          K         K   "       V   '    f�E     �  L  M  f              �  L  N  g              if iteration >= 05��    L                     �%              	       �    L                    �%                     �    L                    �%                     �    L                    �%                     �    L                	   �%             	       �    L         	          �%      	              �    L                   �%                    5�_�  2  4          3  M       ����                                                                                                                                                                                                                                                                                                                i          O         Q                 f�S     �  L  N  g      0        if iteration >= 0 or iteration < 64 then    5��    L                    �%                     �    L                    �%                     �    L                	   �%             	       �    L         	          �%      	              �    L                   �%                    �    L  ,                 �%                    �    L  ,                 �%                    �    L  ,                 �%                    �    L  0                 �%              	       �    M                    �%                    �    M                     �%                     5�_�  3  5          4  O       ����                                                                                                                                                                                                                                                                                                                i          O         Q                 f�h     �  N  P  h                  -- Update kpw�  O  R  h      ,            current_k <= k_const(iteration);   /            current_w <= w_vec(511 downto 480);5��    N                    �%                     �    O                    &                     �    P                    @&                     5�_�  4  6          5  Q       ����                                                                                                                                                                                                                                                                                                                i          Q         O          V       f�j   � �  Q  R  h                  �  Q  S  i              end if;5��    Q                     h&                     �    Q                   p&                    �    Q                   u&                    5�_�  5  7          6  O       ����                                                                                                                                                                                                                                                                                                                i          O         O          V       f��     �  N  R        5��    N                     �%      w               5�_�  6  8          7  A       ����                                                                                                                                                                                                                                                                                                                i          R         R          V       f��     �  A  B  f    �  A  B  f                  -- Update kpw   ,            current_k <= k_const(iteration);   /            current_w <= w_vec(511 downto 480);5��    A                     �$              w       5�_�  7  9          8  B       ����                                                                                                                                                                                                                                                                                                                i          S         Q          V       f��     �  A  B  i       5��    A                     �$                     �    A                     �$                     5�_�  8  :          9  Q       ����                                                                                                                                                                                                                                                                                                                i          Q         Q          V       f��     �  P  T        5��    P                     7&      B               5�_�  9  ;          :  Q        ����                                                                                                                                                                                                                                                                                                                i          Q         Q          V       f��   � �  P  R        5��    P                     7&                     5�_�  :  <          ;  E        ����                                                                                                                                                                                                                                                                                                                i          P         P          V       f��     �  D  F        5��    D                     %      0               5�_�  ;              <  M        ����                                                                                                                                                                                                                                                                                                                i          Q         Q          V       f��   � �  M  N  e    �  M  N  e      /            current_w <= w_vec(511 downto 480);5��    M                     �%              0       5�_�  $          &  %  Q       ����                                                                                                                                                                                                                                                                                                                i                                            f��     �  Q  R  h    �  P  Q  h      /            current_w <= w_vec(511 downto 480);5��    P                     }&              0       5�_�  
                 )    ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f�2     �      d      @    h_register: reg32 port map (rst, clk, enable h7, hv, h_reg);5��      )                  [                      �      +                  ]                      �      *                 \                     �      ,                  ^                      �      +                  ]                      �      *                 \                     �      *                 \                     �      *                 \                     5�_�  �          �  �   p       ����                                                                                                                                                                                                                                                                                                                i             +         +          +    f~P     �   p   q  ^              �   p   r  _              5��    p                      E	                     �    p                  
   E	             
       �    p   	                  N	                     �    p                     M	                     5�_�  �          �  �  
        ����                                                                                                                                                                                                                                                                                                                f             %         9       v   9    fv�     �  
    Y       5��    
                     h                     �    
                     h                     5�_�  �      �  �  �   �   *    ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    ft�   v �   �   �  [      +    signal w_vec: bit_vector(511 downto 0);5��    �   *                  �                     5�_�  �  �      �  �   �   .    ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fs-     �   �   �  [      5    signal current_w: bit_vector(31 downto 0) := msgi5��    �   -                 4                    �    �   2                  9                     �    �   1                 8                    �    �   1                 8                    �    �   1                 8                    5�_�  �  �          �   �   5    ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fs7     �   �   �  [      7    signal current_w: bit_vector(31 downto 0) := msgi()5��    �   5                  <                     5�_�  �  �          �   �   6    ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fs8     �   �   �  [      E    signal current_w: bit_vector(31 downto 0) := msgi(511 downto 480)5��    �   6                  =                     �    �   :                 A                    �    �   :                 A                    �    �   :              
   A             
       5�_�  �  �          �   �   E    ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fs=     �   �   �  [      F    signal current_w: bit_vector(31 downto 0) := msgi(511 downto 480);5��    �   E                  L                     5�_�  �              �  C       ����                                                                                                                                                                                                                                                                                                                f                             V       fsI   t �  B  D        5��    B                     �$      0               5�_�  �          �  �   �       ����                                                                                                                                                                                                                                                                                                                f             '                V   Z    fr[     �   �   �  Y           signal k_const, aux_signals;5��    �                     u                     5�_�  �          �  �   1       ����                                                                                                                                                                                                                                                                                                                g           E   (       E          v       f�     �   0   2        5��    0                      �      !               5�_�  �      �  �  �         ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f��     �            5��                         �      (               5�_�  �          �  �  P       ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f��     �  O  Q  n      !            if iteration  63 then5��    O                    &                     5�_�  X          Z  Y     8    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f��     �      e          �      f              5��                         |                     �                        �                     �                        �                     �                       �                     �                         �                     5�_�  R          T  S   �   $    ����                                                                                                                                                                                                                                                                                                                g           �   :       �   $          $    f�d     �   �   �  e      U    signal op1, op2, op3, op4, op5, op2, op2, op3, op4, op5: bit_vector(31 downto 0);5��    �   &                 z                    5�_�  6  8      9  7     
    ����                                                                                                                                                                                                                                                                                                                g             	         	              f�A     �            5��                         ;      -               5�_�  7              8     
    ����                                                                                                                                                                                                                                                                                                                g             	         	              f�B     �      d    �      d      ,    int2: sigma0 port map(w_vec(i-15), op2);5��                                       -       5�_�  3          5  4         ����                                                                                                                                                                                                                                                                                                                g             	         	              f�,     �      e    �      e      1    int3: adder32 port map(op3, w_vec(i-7), op3);5��                         �              2       5�_�                 �       ����                                                                                                                                                                                                                                                                                                                g           w           w   (       V       f�5     �   �   �  m       5��    �                      A                     �    �                      A                     5�_�  �          �  �  )       ����                                                                                                                                                                                                                                                                                                                H                    E          V       f��     �  (  *  E                  elsif  = 63 then5��    (         	           �"      	               5�_�  W  Y      �  X   �       ����                                                                                                                                                                                                                                                                                                                H           �   +         +          +    f��     �   �   �  4      ,    signal a: bit_vector(31 downto 0) := h0;   /    signal b_in: bit_vector(31 downto 0) := h1;   /    signal c_in: bit_vector(31 downto 0) := h2;   /    signal d_in: bit_vector(31 downto 0) := h3;   /    signal e_in: bit_vector(31 downto 0) := h4;   /    signal f_in: bit_vector(31 downto 0) := h5;   /    signal g_in: bit_vector(31 downto 0) := h6;   /    signal h_in: bit_vector(31 downto 0) := h7;�   �   �  4      /    signal a_in: bit_vector(31 downto 0) := h0;5��    �                     |                     �    �                     �                     �    �                     �                     �    �                                          �    �                     0                     �    �                     ]                     �    �                     �                     �    �                     �                     �    �                     |                     �    �                     �                     �    �                     �                     �    �                                          �    �                     <                     �    �                     l                     �    �                     �                     �    �                     �                     5�_�  X  Z          Y   �   +    ����                                                                                                                                                                                                                                                                                                                H           �   +         +          +    f��     �   �    4      4    a_register: reg32 port map (rst, clk, a, a_reg);   7    b_register: reg32 port map (rst, clk, b_in, b_reg);   7    c_register: reg32 port map (rst, clk, c_in, c_reg);   7    d_register: reg32 port map (rst, clk, d_in, d_reg);   7    e_register: reg32 port map (rst, clk, e_in, e_reg);   7    f_register: reg32 port map (rst, clk, f_in, f_reg);   7    g_register: reg32 port map (rst, clk, g_in, g_reg);   7    h_register: reg32 port map (rst, clk, h_in, h_reg);�   �   �  4      7    a_register: reg32 port map (rst, clk, a_in, a_reg);5��    �   +                  F                     �    �   +                  {                     �    �   +                  �                     �       +                  �                     �      +                                       �      +                  O                     �      +                  �                     �      +                  �                     �    �   +                  F                     �    �   +                  ~                     �    �   +                  �                     �       +                  �                     �      +                  &                     �      +                  ^                     �      +                  �                     �      +                  �                     5�_�  Y  [          Z     !    ����                                                                                                                                                                                                                                                                                                                H                   !                 f��     �      4      A    get_hout: adder32 port map (h7, h_reg, haso(255 downto 224));5��      !                 �                     5�_�  Z  \          [         ����                                                                                                                                                                                                                                                                                                                H                   !                 f�     �    "  4              ao => a,           bo => b_in,           co => c_in,           do => d_in,           eo => e_in,           fo => f_in,           go => g_in,           ho => h_in�      4              ao => a_in,5��                        �!                     �                        �!                     �                        �!                     �                        "                     �                        "                     �                        *"                     �                        ;"                     �                         L"                     �                        �!                     �                        �!                     �                        �!                     �                        "                     �                        %"                     �                        9"                     �                        M"                     �                         a"                     5�_�  [  ]          \           ����                                                                                                                                                                                                                                                                                                                H                                    f�   Z �        4      entity out32 is�   	             end entity out32;�                !architecture Behavior of out32 is�   L   N              component out32 is�   �   �          0    signal a_out: bit_vector(31 downto 0) := h0;�   �   �          0    signal b_out: bit_vector(31 downto 0) := h1;�   �   �          0    signal c_out: bit_vector(31 downto 0) := h2;�   �   �          0    signal d_out: bit_vector(31 downto 0) := h3;�   �   �          0    signal e_out: bit_vector(31 downto 0) := h4;�   �   �          0    signal f_out: bit_vector(31 downto 0) := h5;�   �   �          0    signal g_out: bit_vector(31 downto 0) := h6;�   �   �          0    signal h_out: bit_vector(31 downto 0) := h7;�   �   �          7    a_outister: out32 port map (rst, clk, a_in, a_out);�   �             7    b_outister: out32 port map (rst, clk, b_in, b_out);�   �            7    c_outister: out32 port map (rst, clk, c_in, c_out);�               7    d_outister: out32 port map (rst, clk, d_in, d_out);�              7    e_outister: out32 port map (rst, clk, e_in, e_out);�              7    f_outister: out32 port map (rst, clk, f_in, f_out);�              7    g_outister: out32 port map (rst, clk, g_in, g_out);�              7    h_outister: out32 port map (rst, clk, h_in, h_out);�              >    get_aout: adder32 port map (h0, a_out, haso(31 downto 0));�    	          ?    get_bout: adder32 port map (h1, b_out, haso(63 downto 32));�    
          ?    get_cout: adder32 port map (h2, c_out, haso(95 downto 64));�  	            @    get_dout: adder32 port map (h3, d_out, haso(127 downto 96));�  
            A    get_eout: adder32 port map (h4, e_out, haso(159 downto 128));�              A    get_fout: adder32 port map (h5, f_out, haso(191 downto 160));�              A    get_gout: adder32 port map (h6, g_out, haso(223 downto 192));�              A    get_hout: adder32 port map (h7, h_out, haso(255 downto 224));�                      ai => a_out,�                      bi => b_out,�                      ci => c_out,�                      di => d_out,�                      ei => e_out,�                      fi => f_out,�                      gi => g_out,�                      hi => h_out,5��                        0                     �    	                    �                     �                        �                     �    L                    W                    �    �                    �                    �    �                    .                    �    �                    _                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    #                    �    �                    T                    �    �                    !                    �    �                    +                    �    �   2                 M                    �    �                    Y                    �    �                    c                    �    �   2                 �                    �    �                    �                    �    �                    �                    �    �   2                 �                    �                        �                    �                        �                    �       2                 �                    �                                           �                                           �      2                 -                    �                       9                    �                       C                    �      2                 e                    �                       q                    �                       {                    �      2                 �                    �                       �                    �                       �                    �      2                 �                    �      &                                     �      &                 A                    �      &                 �                    �    	  &                 �                    �    
  &                                      �      &                 D                     �      &                 �                     �      &                 �                     �                       !                    �                       '!                    �                       <!                    �                       Q!                    �                       f!                    �                       {!                    �                       �!                    �                       �!                    5�_�  \  ^          ]         ����                                                                                                                                                                                                                                                                                                                H                   !                 f�6     �      4              ai => a_,           bi => b_,           ci => c_,           di => d_,           ei => e_,           fi => f_,           gi => g_,           hi => h_,5��                        !                     �                        $!                     �                        6!                     �                        H!                     �                        Z!                     �                        l!                     �                        ~!                     �                        �!                     5�_�  ]  _          ^         ����                                                                                                                                                                                                                                                                                                                H                                    f�:     �    "  4              ao => a_,           bo => b_,           co => c_,           do => d_,           eo => e_,           fo => f_,           go => g_,           ho => h_�      4    �    #  4   	           ao => a_out,           bo => b_out,           co => c_out,           do => d_out,           eo => e_out,           fo => f_out,           go => g_out,           ho => h_out       );5��                        �!                     �                        �!                     �                        �!                     �                        �!                     �                        "                     �                        "                     �                        *"                     �                         <"                     �                        �!                     �                        �!                     �                        �!                     �                        �!                     �                        "                     �                        '"                     �                        <"                     �                         Q"                     5�_�  ^  `          _         ����                                                                                                                                                                                                                                                                                                                H                                    f�@     �      4              ai => a,           bi => b,           ci => c,           di => d,           ei => e,           fi => f,           gi => g,           hi => h,�      4    �      4   	           ai => ain,           bi => bin,           ci => cin,           di => din,           ei => ein,           fi => fin,           gi => gin,           hi => hin,           kpw => current_kpw,5��                        !                     �                        "!                     �                        3!                     �                        D!                     �                        U!                     �                        f!                     �                        w!                     �                        �!                     �                        !                     �                        $!                     �                        7!                     �                        J!                     �                        ]!                     �                        p!                     �                        �!                     �                        �!                     5�_�  _  a          `         ����                                                                                                                                                                                                                                                                                                                H                                    f�I     �      4              ai => a_in,�      4              bi => b_in,           ci => c_in,           di => d_in,           ei => e_in,           fi => f_in,           gi => g_in,           hi => h_in,5��                        !                     �                        %!                     �                        9!                     �                        M!                     �                        a!                     �                        u!                     �                        �!                     �                        �!                     5�_�  `  b          a  %       ����                                                                                                                                                                                                                                                                                                                H                                    f�X     �  %  &  4              �  %  '  5                  variable i5��    %                     �"                     �    %                    �"                    �    %                     �"                     �    %                    �"              	       �    &                 
   �"              
       5�_�  a  c          b  '       ����                                                                                                                                                                                                                                                                                                                H           �                   V       f�^     �  &  (  6              variable iteration5��    &                    �"                     �    &                   �"                    5�_�  b  d          c         ����                                                                                                                                                                                                                                                                                                                H           �                   V       f�q     �   �    6      :    -- a_outister: out32 port map (rst, clk, a_in, a_out);   :    -- b_outister: out32 port map (rst, clk, b_in, b_out);   :    -- c_outister: out32 port map (rst, clk, c_in, c_out);   :    -- d_outister: out32 port map (rst, clk, d_in, d_out);   :    -- e_outister: out32 port map (rst, clk, e_in, e_out);   :    -- f_outister: out32 port map (rst, clk, f_in, f_out);   :    -- g_outister: out32 port map (rst, clk, g_in, g_out);   :    -- h_outister: out32 port map (rst, clk, h_in, h_out);5��    �                           �      �      5�_�  c  e          d   �       ����                                                                                                                                                                                                                                                                                                                H           �                   V       f�t     �   �   �  6      <    -- counter: counter_6bit port map (clk, rst, iteration);5��    �                     �      :       =       5�_�  d  f          e   �       ����                                                                                                                                                                                                                                                                                                                H           �                   V       f�   [ �   �   �  6              �   �   �  7          -- Registers5��    �                                           �    �                                         �    �                    "                    5�_�  e  g          f  (       ����                                                                                                                                                                                                                                                                                                                H           �                   V       f��     �  '  )  7      $        variable iteration: integer 5��    '                 
   �"              
       5�_�  f  h          g  (   #    ����                                                                                                                                                                                                                                                                                                                H           �                   V       f��     �  (  )  7    �  (  )  7      ,        	variable i : integer range 0 to 64;5��    (                     �"              -       5�_�  g  i          h  )   	    ����                                                                                                                                                                                                                                                                                                                H           �                   V       f��     �  (  *  8      +        variable i : integer range 0 to 64;5��    (                    �"                     5�_�  h  j          i  (       ����                                                                                                                                                                                                                                                                                                                H           �                   V       f��     �  '  )        5��    '                     �"      %               5�_�  i  k          j  (       ����                                                                                                                                                                                                                                                                                                                H           �                   V       f��     �  '  )  7      3        variable iteration : integer range 0 to 64;5��    '                    �"                     5�_�  j  l          k  (       ����                                                                                                                                                                                                                                                                                                                H           �                   V       f��     �  '  )        5��    '                     �"      4               5�_�  k  m          l  &        ����                                                                                                                                                                                                                                                                                                                H           �                   V       f��     �  &  '  6    �  %  &  6      3        variable iteration : integer range 0 to 64;5��    %                     �"              4       5�_�  l  n          m  &       ����                                                                                                                                                                                                                                                                                                                H           �                   V       f��     �  %  '  7      /    variable iteration : integer range 0 to 64;5��    %                    �"                     5�_�  m  o          n  &       ����                                                                                                                                                                                                                                                                                                                H          *          4           V        f��     �  %  '  7      3        variable iteration : integer range 0 to 64;5��    %                    �"                     5�_�  n  p          o  *        ����                                                                                                                                                                                                                                                                                                                H          P         *                 f��     �  )  5        �  *  +  ,    �  )  *  ,   '   '            	if (rising_edge(clk)) then   '                    if (rst = '1') then                           i := 0;   $                        done <= '0';                       end if;       1                    if (rst = '0' and i = 0) then   +                        ain <= x"6a09e667";   +                        bin <= x"bb67ae85";   +                        cin <= x"3c6ef372";   +                        din <= x"a54ff53a";   2                        ein <= x"510e527f";          +                        fin <= x"9b05688c";   +                        gin <= x"1f83d9ab";   +                        hin <= x"5be0cd19";   (                        kpwin <= KPW(0);                       end if;       /                    if (i /= 0 and i < 64) then   $                        ain <= aout;   $                        bin <= bout;   $                        cin <= cout;   $                        din <= dout;   $                        ein <= eout;   $                        fin <= fout;   $                        gin <= gout;   $                        hin <= hout;   (                        kpwin <= KPW(i);                       end if;       $                    if (i = 64) then   $                        done <= '1';                       end if;                          2                    if (rst = '0' and i < 64) then                        	i := i + 1;                       end if;                   end if;           end process; 5��    )                     �"                    �    )              '       �"              H      5�_�  o  q          p  *       ����                                                                                                                                                                                                                                                                                                                H          P         *                 f��     �  )  +  S          	if (rising_edge(clk)) then5��    )                     �"                     5�_�  p  r          q  )        ����                                                                                                                                                                                                                                                                                                                H          O         )                 f��     �  (  *        5��    (                     �"                     5�_�  q  s          r  )       ����                                                                                                                                                                                                                                                                                                                H          O         )                 f��     �  (  *  R          if (rising_edge(clk)) then5��    (                    �"                     5�_�  r  t          s  *       ����                                                                                                                                                                                                                                                                                                                H          O         )                 f��     �  )  +  R              if (rst = '1') then5��    )                    #                     5�_�  s  u          t  +       ����                                                                                                                                                                                                                                                                                                                H          O         )                 f��     �  *  ,  R                  i := 0;5��    *                    ;#                     �    *                    :#                     �    *                    9#                     �    *                    8#                     �    *                    7#                     �    *                    6#                     �    *                    5#                     �    *                    4#                     �    *                    3#                     �    *                    2#                     �    *                    1#                     �    *                    0#                     5�_�  t  v          u  +       ����                                                                                                                                                                                                                                                                                                                H          O         )                 f��     �  *  ,  R                  iteration := 0;5��    *                    1#                     5�_�  u  w          v  ,       ����                                                                                                                                                                                                                                                                                                                H          O         )                 f��     �  +  -  R                  done <= '0';5��    +                    L#                     5�_�  v  x          w  -       ����                                                                                                                                                                                                                                                                                                                H          O         )                 f��     �  ,  .  R              end if;5��    ,                    a#                     5�_�  w  y          x  /       ����                                                                                                                                                                                                                                                                                                                H          O         )                 f��     �  .  0  R      %        if (rst = '0' and i = 0) then5��    .                   n#                    5�_�  x  z          y  0       ����                                                                                                                                                                                                                                                                                                                H          1         8                 f��     �  /  1  R                  ain <= x"6a09e667";5��    /                    �#                     �    /                    �#                     �    /                    �#                     �    /                    �#                     �    /                    �#                     �    /                    �#                     �    /                    �#                     �    /                    �#                     �    /                    �#                     �    /                    �#                     �    /                    �#                     �    /                    �#                     5�_�  y  {          z  1       ����                                                                                                                                                                                                                                                                                                                H          1         8                 f��     �  0  2  R                  bin <= x"bb67ae85";5��    0                    �#                     �    0                    �#                     �    0                    �#                     �    0                    �#                     �    0                    �#                     �    0                    �#                     �    0                    �#                     �    0                    �#                     �    0                    �#                     �    0                    �#                     �    0                    �#                     �    0                    �#                     5�_�  z  |          {  2       ����                                                                                                                                                                                                                                                                                                                H          1         8                 f��     �  1  3  R                  cin <= x"3c6ef372";5��    1                    �#                     �    1                    �#                     �    1                    �#                     �    1                    �#                     �    1                    �#                     �    1                    �#                     �    1                    �#                     �    1                    �#                     �    1                    �#                     �    1                    �#                     �    1                    �#                     �    1                    �#                     5�_�  {  }          |  3       ����                                                                                                                                                                                                                                                                                                                H          1         8                 f��     �  2  4  R                  din <= x"a54ff53a";5��    2                    $                     �    2                    $                     �    2                    $                     �    2                    $                     �    2                    $                     �    2                    $                     �    2                    $                     �    2                     $                     �    2                    �#                     �    2                    �#                     �    2                    �#                     �    2                    �#                     5�_�  |  ~          }  4       ����                                                                                                                                                                                                                                                                                                                H          1         8                 f��     �  3  5  R      &            ein <= x"510e527f";       5��    3                    '$                     �    3                    &$                     �    3                    %$                     �    3                    $$                     �    3                    #$                     �    3                    "$                     �    3                    !$                     �    3                     $                     �    3                    $                     �    3                    $                     �    3                    $                     �    3                    $                     5�_�  }            ~  5       ����                                                                                                                                                                                                                                                                                                                H          1         8                 f��     �  4  6  R                  fin <= x"9b05688c";5��    4                    N$                     �    4                    M$                     �    4                    L$                     �    4                    K$                     �    4                    J$                     �    4                    I$                     �    4                    H$                     �    4                    G$                     �    4                    F$                     �    4                    E$                     �    4                    D$                     �    4                    C$                     5�_�  ~  �            6       ����                                                                                                                                                                                                                                                                                                                H          1         8                 f��     �  5  7  R                  gin <= x"1f83d9ab";5��    5                    n$                     �    5                    m$                     �    5                    l$                     �    5                    k$                     �    5                    j$                     �    5                    i$                     �    5                    h$                     �    5                    g$                     �    5                    f$                     �    5                    e$                     �    5                    d$                     �    5                    c$                     5�_�    �          �  7       ����                                                                                                                                                                                                                                                                                                                H          1         8                 f�      �  6  8  R                  hin <= x"5be0cd19";5��    6                    �$                     �    6                    �$                     �    6                    �$                     �    6                    �$                     �    6                    �$                     �    6                    �$                     �    6                    �$                     �    6                    �$                     �    6                    �$                     �    6                    �$                     �    6                    �$                     �    6                    �$                     5�_�  �  �          �  8       ����                                                                                                                                                                                                                                                                                                                H          0         7                 f�     �  7  9  R                  kpwin <= KPW(0);5��    7                    �$                     �    7                    �$                     �    7                    �$                     �    7                    �$                     �    7                    �$                     �    7                    �$                     �    7                    �$                     �    7                    �$                     �    7                    �$                     �    7                    �$                     �    7                    �$                     �    7                    �$                     5�_�  �  �          �  0       ����                                                                                                                                                                                                                                                                                                                H          1         7                 f�	     �  /  8  R                  ain <= ;               bin <= h0;               cin <= h0;               din <= h0;               ein <= h0;                      fin <= h0;               gin <= h0;               hin <= h0;�  /  1  R                  ain <= h0;5��    /                    �#                     �    0                    �#                     �    1                    �#                     �    2                    �#                     �    3                    �#                     �    4                    $                     �    5                    ($                     �    6                    =$                     �    /                    �#                     �    0                    �#                     �    1                    �#                     �    2                    �#                     �    3                    �#                     �    4                    $                     �    5                    4$                     �    6                    K$                     5�_�  �  �          �  1       ����                                                                                                                                                                                                                                                                                                                H          0         7                 f�     �  0  8  R                  bin <= h1;               cin <= h2;               din <= h3;               ein <= h4;                      fin <= h5;               gin <= h6;               hin <= h7;5��    0                   �#                    �    1                   �#                    �    2                   �#                    �    3                    $                    �    4                   $                    �    5                   5$                    �    6                   L$                    5�_�  �  �          �  0       ����                                                                                                                                                                                                                                                                                                                H          0         7                 f�     �  /  1  R                  a_in <= h0;�  0  8  R                  b_in <= h1;               c_in <= h2;               d_in <= h3;               e_in <= h4;                      f_in <= h5;               g_in <= h6;               h_in <= h7;5��    /                    �#                     �    0                    �#                     �    1                    �#                     �    2                    �#                     �    3                    �#                     �    4                    $                     �    5                    4$                     �    6                    L$                     5�_�  �  �          �  8       ����                                                                                                                                                                                                                                                                                                                H          0         7                 f�     �  7  9  R      "            current_kpw <= KPW(0);5��    7                   c$                    �    7                    f$                     �    7                    e$                     �    7                    d$                     �    7                   c$                    �    7                   c$                    �    7                   c$                    5�_�  �  �          �  8       ����                                                                                                                                                                                                                                                                                                                H          0         7                 f�     �  7  9  R      &            current_kpw <= kpw_vec(0);5��    7                   r$                    �    7                    t$                     �    7                    s$                     �    7                   r$                    �    7                   r$                    �    7                   r$                    5�_�  �  �          �  /       ����                                                                                                                                                                                                                                                                                                                H          0         7                 f�#     �  .  0  R      -        if (rst = '0' and iteration = 0) then5��    .                   �#                    �    .                    �#                     �    .                	   �#             	       �    .         	          �#      	              �    .                	   �#             	       5�_�  �  �          �  9       ����                                                                                                                                                                                                                                                                                                                H          0         7                 f�'     �  8  :  R              end if;5��    8                    �$                     5�_�  �  �          �  ;       ����                                                                                                                                                                                                                                                                                                                H          ;         ;          V       f�)     �  :  <  R      #        if (i /= 0 and i < 64) then5��    :                    �$                     5�_�  �  �          �  ;        ����                                                                                                                                                                                                                                                                                                                H          ;         ;          V       f�6     �  :  <  R      ;        iterationf (iteration /= 0 and iteration < 64) then5��    :                	   �$             	       �    :                	   �$             	       �    :  '              	   �$             	       5�_�  �  �          �  ;       ����                                                                                                                                                                                                                                                                                                                H          <         D                 f�7     �  :  <  R      3        if (iteration /= 0 and iteration < 64) then5��    :         
          �$      
              5�_�  �  �          �  <       ����                                                                                                                                                                                                                                                                                                                H          <         D                 f�@     �  ;  =  R                  ain <= aout;5��    ;                    �$                     �    ;                    �$                     �    ;                    �$                     �    ;                    �$                     �    ;                    �$                     �    ;                    �$                     �    ;                    �$                     �    ;                    �$                     �    ;                    �$                     �    ;                    �$                     �    ;                    �$                     �    ;                    �$                     5�_�  �  �          �  =       ����                                                                                                                                                                                                                                                                                                                H          <         D                 f�C     �  <  >  R                  bin <= bout;5��    <                    �$                     �    <                    �$                     �    <                    �$                     �    <                    �$                     �    <                    �$                     �    <                    �$                     �    <                    �$                     �    <                    �$                     �    <                    �$                     �    <                    �$                     �    <                    �$                     �    <                    �$                     5�_�  �  �          �  >       ����                                                                                                                                                                                                                                                                                                                H          <         D                 f�D     �  =  ?  R                  cin <= cout;5��    =                    %                     �    =                    %                     �    =                    %                     �    =                    %                     �    =                    %                     �    =                    %                     �    =                    %                     �    =                    %                     �    =                    %                     �    =                    %                     �    =                    
%                     �    =                    	%                     5�_�  �  �          �  ?       ����                                                                                                                                                                                                                                                                                                                H          <         D                 f�E     �  >  @  R                  din <= dout;5��    >                    -%                     �    >                    ,%                     �    >                    +%                     �    >                    *%                     �    >                    )%                     �    >                    (%                     �    >                    '%                     �    >                    &%                     �    >                    %%                     �    >                    $%                     �    >                    #%                     �    >                    "%                     5�_�  �  �          �  @       ����                                                                                                                                                                                                                                                                                                                H          <         D                 f�F     �  ?  A  R                  ein <= eout;5��    ?                    F%                     �    ?                    E%                     �    ?                    D%                     �    ?                    C%                     �    ?                    B%                     �    ?                    A%                     �    ?                    @%                     �    ?                    ?%                     �    ?                    >%                     �    ?                    =%                     �    ?                    <%                     �    ?                    ;%                     5�_�  �  �          �  A       ����                                                                                                                                                                                                                                                                                                                H          <         D                 f�G     �  @  B  R                  fin <= fout;5��    @                    _%                     �    @                    ^%                     �    @                    ]%                     �    @                    \%                     �    @                    [%                     �    @                    Z%                     �    @                    Y%                     �    @                    X%                     �    @                    W%                     �    @                    V%                     �    @                    U%                     �    @                    T%                     5�_�  �  �          �  B       ����                                                                                                                                                                                                                                                                                                                H          <         D                 f�I     �  A  C  R                  gin <= gout;5��    A                    x%                     �    A                    w%                     �    A                    v%                     �    A                    u%                     �    A                    t%                     �    A                    s%                     �    A                    r%                     �    A                    q%                     �    A                    p%                     �    A                    o%                     �    A                    n%                     �    A                    m%                     5�_�  �  �          �  C       ����                                                                                                                                                                                                                                                                                                                H          <         D                 f�J     �  B  D  R                  hin <= hout;5��    B                    �%                     �    B                    �%                     �    B                    �%                     �    B                    �%                     �    B                    �%                     �    B                    �%                     �    B                    �%                     �    B                    �%                     �    B                    �%                     �    B                    �%                     �    B                    �%                     �    B                    �%                     5�_�  �  �          �  D       ����                                                                                                                                                                                                                                                                                                                H          <         D                 f�K     �  C  E  R                  kpwin <= KPW(i);5��    C                    �%                     �    C                    �%                     �    C                    �%                     �    C                    �%                     �    C                    �%                     �    C                    �%                     �    C                    �%                     �    C                    �%                     �    C                    �%                     �    C                    �%                     �    C                    �%                     �    C                    �%                     5�_�  �  �          �  E       ����                                                                                                                                                                                                                                                                                                                H          <         C                 f�L     �  D  F  R              end if;5��    D                    �%                     5�_�  �  �          �  <       ����                                                                                                                                                                                                                                                                                                                H          <         C                 f�T     �  ;  =  R                  a_in <= aout;�  <  D  R                  b_in <= bout;               c_in <= cout;               d_in <= dout;               e_in <= eout;               f_in <= fout;               g_in <= gout;               h_in <= hout;5��    ;                    �$                     �    <                    �$                     �    =                    %                     �    >                    &%                     �    ?                    @%                     �    @                    Z%                     �    A                    t%                     �    B                    �%                     5�_�  �  �          �  <       ����                                                                                                                                                                                                                                                                                                                H          <         C                 f�X     �  ;  =  R                  a_in <= a_out;�  <  D  R                  b_in <= b_out;               c_in <= c_out;               d_in <= d_out;               e_in <= e_out;               f_in <= f_out;               g_in <= g_out;               h_in <= h_out;5��    ;                    �$                     �    <                    �$                     �    =                    %                     �    >                    1%                     �    ?                    L%                     �    @                    g%                     �    A                    �%                     �    B                    �%                     5�_�  �  �          �  D       ����                                                                                                                                                                                                                                                                                                                H          <         C                 f�[     �  C  E  R                   kpwin <= kpw_vec(i);5��    C                   �%                    �    C                    �%                     �    C                    �%                     �    C                   �%                    �    C                   �%                    �    C                   �%                    5�_�  �  �          �  D       ����                                                                                                                                                                                                                                                                                                                H          <         C                 f�^     �  C  E  R      &            current_kpw <= kpw_vec(i);5��    C                   �%                    �    C                    �%                     �    C                    �%                     �    C                   �%                    �    C                   �%                    �    C                   �%                    5�_�  �  �          �  D   #    ����                                                                                                                                                                                                                                                                                                                H          <         C                 f�a     �  C  E  R      .            current_kpw <= kpw_vec(iteration);5��    C  #                 �%                    �    C  %                  �%                     �    C  $                  �%                     �    C  #              	   �%             	       �    C  #       	          �%      	              �    C  #              	   �%             	       5�_�  �  �          �  G       ����                                                                                                                                                                                                                                                                                                                H          <         C                 f�d     �  F  H  R              if (i = 64) then5��    F                    �%                     5�_�  �  �          �  H       ����                                                                                                                                                                                                                                                                                                               H         <         C                 f�f     �  G  I  R                  done <= '1';5��    G                    &                     5�_�  �      �      �  H       ����                                                                                                                                                                                                                                                                                                               H         <         C                 f�f     �  G  J  R                   done <= '1'; end if;5��    G                  &                    5�_�  �  �      �  �  I       ����                                                                                                                                                                                                                                                                                                               H         <         C                 f�h     �  H  J  R              end if;5��    H                    &                     5�_�  �  �          �  K       ����                                                                                                                                                                                                                                                                                                               H         <         C                 f�k     �  J  L  R      &        if (rst = '0' and i < 64) then5��    J                    B&                     5�_�  �  �          �  L       ����                                                                                                                                                                                                                                                                                                               H         <         C                 f�l     �  K  M  R                  i := i + 1;5��    K                    u&                     �    K                    t&                     �    K                    s&                     �    K                    r&                     �    K                    q&                     �    K                    p&                     �    K                    o&                     �    K                    n&                     �    K                    m&                     5�_�  �  �          �  M       ����                                                                                                                                                                                                                                                                                                               H         <         C                 f�m     �  L  N  R              end if;5��    L                    �&                     5�_�  �  �          �  N       ����                                                                                                                                                                                                                                                                                                               H         <         C                 f�p     �  M  O  R          end if;5��    M                    �&                     5�_�  �  �          �  O       ����                                                                                                                                                                                                                                                                                                               H         <         C                 f�q     �  N  P  R          end process; 5��    N                    �&                    5�_�  �  �          �  O       ����                                                                                                                                                                                                                                                                                                               H         <         C                 f�w     �  N  P  R      end process; 5��    N                     �&                     5�_�  �  �          �  L       ����                                                                                                                                                                                                                                                                                                               H         <         C                 f�{     �  K  M  R                  iteration := i + 1;5��    K                   m&                    �    K                    o&                     �    K                    n&                     �    K                	   m&             	       �    K         	          m&      	              �    K                	   m&             	       5�_�  �  �          �  L       ����                                                                                                                                                                                                                                                                                                               H         <         C                 f�~     �  K  M  R      '            iteration := iteration + 1;5��    K                   z&                    �    K                    |&                     �    K                    {&                     �    K                	   z&             	       �    K         	          z&      	              �    K                	   z&             	       5�_�  �  �          �  K       ����                                                                                                                                                                                                                                                                                                               H         <         C                 f��     �  J  L  R      .        if (rst = '0' and iteration < 64) then5��    J                   T&                    �    J                    V&                     �    J                    U&                     �    J                	   T&             	       �    J         	          T&      	              �    J                	   T&             	       5�_�  �  �          �  G       ����                                                                                                                                                                                                                                                                                                               H         <         C                 f��   \ �  F  H  R               if (iteration = 64) then5��    F                   �%                    �    F                    �%                     �    F                    �%                     �    F                	   �%             	       �    F         	          �%      	              �    F                	   �%             	       5�_�  �  �          �   M        ����                                                                                                                                                                                                                                                                                                               @         4         ;                 f��     �   L   U        5��    L                      I      �               5�_�  �  �          �   M        ����                                                                                                                                                                                                                                                                                                               9          6                     V       f��     �   L   T        5��    L                      I      �               5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                              V       f��   ] �       7        5��            6                       8              5�_�  �  �          �   ;       ����                                                                                                                                                                                                                                                                                                                                              V       f��   ^ �   :   <        5��    :                            $               5�_�  �  �          �   ;       ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   :   <        1    signal a_in, : bit_vector(31 downto 0) := h0;5��    :                     �                     5�_�  �  �          �   ;       ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   ;   <      �   :   <        7    signal a_in, a_in, : bit_vector(31 downto 0) := h0;5��    :                     �                     5�_�  �  �          �   ;       ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   ;   <      �   :   <        =    signal a_in, a_in, a_in, : bit_vector(31 downto 0) := h0;5��    :                     �                     5�_�  �  �          �   ;       ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   ;   <      �   :   <        C    signal a_in, a_in, a_in, a_in, : bit_vector(31 downto 0) := h0;5��    :                     �                     5�_�  �  �          �   ;   "    ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   ;   <      �   :   <        I    signal a_in, a_in, a_in, a_in, a_in, : bit_vector(31 downto 0) := h0;5��    :   #                  �                     5�_�  �  �          �   ;   (    ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   ;   <      �   :   <        O    signal a_in, a_in, a_in, a_in, a_in, a_in, : bit_vector(31 downto 0) := h0;5��    :   )                  �                     5�_�  �  �          �   ;   .    ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   ;   <      �   :   <        U    signal a_in, a_in, a_in, a_in, a_in, a_in, a_in, : bit_vector(31 downto 0) := h0;5��    :   /                  �                     5�_�  �  �          �   ;   4    ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   ;   <      �   :   <        [    signal a_in, a_in, a_in, a_in, a_in, a_in, a_in, a_in, : bit_vector(31 downto 0) := h0;5��    :   5                  �                     5�_�  �  �          �   ;   :    ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   ;   <      �   :   <        a    signal a_in, a_in, a_in, a_in, a_in, a_in, a_in, a_in, a_in, : bit_vector(31 downto 0) := h0;5��    :   ;                  �                     5�_�  �  �          �   ;   @    ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   :   <        `    signal a_in, a_in, a_in, a_in, a_in, a_in, a_in, a_in, a_in,: bit_vector(31 downto 0) := h0;5��    :   @                  �                     5�_�  �  �          �   ;   ?    ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   :   <        _    signal a_in, a_in, a_in, a_in, a_in, a_in, a_in, a_in, a_in: bit_vector(31 downto 0) := h0;5��    :   ?                  �                     5�_�  �  �          �   ;       ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   :   <        _    signal a_in, b_in, a_in, a_in, a_in, a_in, a_in, a_in, a_in: bit_vector(31 downto 0) := h0;5��    :                    �                    5�_�  �  �          �   ;       ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   :   <        _    signal a_in, b_in, c_in, a_in, a_in, a_in, a_in, a_in, a_in: bit_vector(31 downto 0) := h0;5��    :                    �                    5�_�  �  �          �   ;       ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   :   <        _    signal a_in, b_in, c_in, d_in, a_in, a_in, a_in, a_in, a_in: bit_vector(31 downto 0) := h0;5��    :                    �                    5�_�  �  �          �   ;   #    ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   :   <        _    signal a_in, b_in, c_in, d_in, e_in, a_in, a_in, a_in, a_in: bit_vector(31 downto 0) := h0;5��    :   #                 �                    5�_�  �  �          �   ;   )    ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   :   <        _    signal a_in, b_in, c_in, d_in, e_in, f_in, a_in, a_in, a_in: bit_vector(31 downto 0) := h0;5��    :   )                 �                    5�_�  �  �          �   ;   /    ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   :   <        _    signal a_in, b_in, c_in, d_in, e_in, f_in, g_in, a_in, a_in: bit_vector(31 downto 0) := h0;5��    :   /                 �                    5�_�  �  �          �   ;   5    ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f��     �   :   <        _    signal a_in, b_in, c_in, d_in, e_in, f_in, g_in, h_in, a_in: bit_vector(31 downto 0) := h0;5��    :   5                 �                    5�_�  �  �          �   ;   ;    ����                                                                                                                                                                                                                                                                                                                         ;          ;          v       f�     �   :   <        [    signal a_in, b_in, c_in, d_in, e_in, f_in, g_in, h_in, : bit_vector(31 downto 0) := h0;5��    :   ;                  �                     5�_�  �  �          �   ;   9    ����                                                                                                                                                                                                                                                                                                                         <   .       B   /       V   9    f�	     �   :   <        Y    signal a_in, b_in, c_in, d_in, e_in, f_in, g_in, h_in: bit_vector(31 downto 0) := h0;5��    :   9                  �                     5�_�  �  �          �   <        ����                                                                                                                                                                                                                                                                                                                �          <   .       <   /       V   9    f�     �   ;   C        5��    ;                      �      P              5�_�  �  �          �   ;   /    ����                                                                                                                                                                                                                                                                                                                �          <          <          V       f�'     �   ;   <      �   ;   <        Y    signal a_in, b_in, c_in, d_in, e_in, f_in, g_in, h_in: bit_vector(31 downto 0) := h0;5��    ;                      �              Z       5�_�  �  �  �      �   <        ����                                                                                                                                                                                                                                                                                                                �          <          <          V       f�.     �   ;   =        a    signal a_out, b_out, c_out, d_out, e_out, f_out, g_out, h_out: bit_vector(31 downto 0) := h0;5��    ;                    �                    �    ;                    �                    �    ;                    �                    �    ;   "                 �                    �    ;   )                                     �    ;   0                 	                    �    ;   7                                     �    ;   >                                     5�_�  �  �          �   =       ����                                                                                                                                                                                                                                                                                                                �          �          �          V       f�0   _ �   <   E        5��    <                      ;      �              5�_�  �  �  �      �   �        ����                                                                                                                                                                                                                                                                                                                �          �          �          V       f�X     �   �   �        �   �   �          entity somador32 is   
    port (   '        a : in bit_vector(31 downto 0);   '        b : in bit_vector(31 downto 0);   '        r : out bit_vector(31 downto 0)       );   end entity somador32;       'architecture behavioral of somador32 is   +    signal carry : bit_vector(31 downto 0);   begin   "    sum: for i in 0 to 30 generate   +        r(i) <= A(i) xor B(i) xor carry(i);   T        carry(i+1) <= (A(i) and B(i)) or (A(i) and carry(i)) or (B(i) and carry(i));       end generate;       +    r(31) <= A(31) xor B(31) xor carry(31);          end architecture behavioral;    5��    �                      �                    5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                �          �          �          V       f�b   ` �                  component somador32  is�   �   �          9        	make3: somador32 port map(op3, w_vec(i-7), op3);�   �   �          2        	make4: somador32 port map(op3, op2, op4);�   �   �          :        	make5: somador32 port map(op4, w_vec(i-16), op5);�   �   �          2        	make1: somador32 port map(op1, op2, op3);�   �   �          @    get_aout: somador32 port map (h0, a_out, haso(31 downto 0));�   �   �          A    get_bout: somador32 port map (h1, b_out, haso(63 downto 32));�   �   �          A    get_cout: somador32 port map (h2, c_out, haso(95 downto 64));�   �   �          B    get_dout: somador32 port map (h3, d_out, haso(127 downto 96));�   �   �          C    get_eout: somador32 port map (h4, e_out, haso(159 downto 128));�   �   �          C    get_fout: somador32 port map (h5, f_out, haso(191 downto 160));�   �   �          C    get_gout: somador32 port map (h6, g_out, haso(223 downto 192));�   �   �          C    get_hout: somador32 port map (h7, h_out, haso(255 downto 224));5��                     	                	       �    �                 	   �             	       �    �                 	                	       �    �                 	   K             	       �    �                 	   W             	       �    �                 	   �             	       �    �                 	   $             	       �    �                 	   f             	       �    �                 	   �             	       �    �                 	   �             	       �    �                 	   /             	       �    �                 	   s             	       �    �                 	   �             	       5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                �          �          �          V       f�r     �   �   �        5��    �                      �      '              5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                �          �          �          V       f�s   a �   �   �        5��    �                      �                     5�_�  �  �          �   ;   R    ����                                                                                                                                                                                                                                                                                                                �          �          �          V       f�P     �   :   <        S    signal a_in, b_in, c_in, d_in, e_in, f_in, g_in, h_in: bit_vector(31 downto 0);5��    :   R                  �                     5�_�  �  �          �   <   Z    ����                                                                                                                                                                                                                                                                                                                �          �                     V        f�T   b �   ;   =        [    signal a_out, b_out, c_out, d_out, e_out, f_out, g_out, h_out: bit_vector(31 downto 0);5��    ;   Z                  /                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                �          �                     V        f�R     �   �   �        entity somador is5��    �                     �                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                �          �                     V        f�V     �   �   �        end entity somador;5��    �                     7                     �    �                     6                     5�_�  �  �          �   �   $    ����                                                                                                                                                                                                                                                                                                                �          �                     V        f�X   c �   �   �        %architecture behavioral of somador is5��    �   #                  \                     �    �   "                  [                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                �          �                     V        f�]     �                  component somadoris5��                         &                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                �          �          �                 f�^     �                  component somador is5��                         &                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                �          �          �                 f�f     �   �   �        7        	make3: somador port map(op3, w_vec(i-7), op3);   0        	make4: somador port map(op3, op2, op4);   8        	make5: somador port map(op4, w_vec(i-16), op5);5��    �                     �                     �    �                                          �    �                     ?                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                �          �          �                 f�i     �   �   �        1        	make1: somador2 port map(op1, op2, op3);5��    �                     I                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                �          �          �                 f�i     �   �   �        0        	make1: somador port map(op1, op2, op3);5��    �                     I                     5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                �                                           f�l   d �   �   �        >    get_aout: somador port map (h0, a_out, haso(31 downto 0));   ?    get_bout: somador port map (h1, b_out, haso(63 downto 32));   ?    get_cout: somador port map (h2, c_out, haso(95 downto 64));   @    get_dout: somador port map (h3, d_out, haso(127 downto 96));   A    get_eout: somador port map (h4, e_out, haso(159 downto 128));   A    get_fout: somador port map (h5, f_out, haso(191 downto 160));   A    get_gout: somador port map (h6, g_out, haso(223 downto 192));   A    get_hout: somador port map (h7, h_out, haso(255 downto 224));5��    �                     �                     �    �                     �                     �    �                     *                     �    �                     j                     �    �                     �                     �    �                     �                     �    �                     /                     �    �                     q                     5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                �                                           f��   e �              entity multisteps_v0 is5��                         :                      �                        <                     5�_�  �              �          ����                                                                                                                                                                                                                                                                                                                �                                           f��   f �   
           end multisteps_v0;5��    
                     �                      5�_�  �          �  �          ����                                                                                                                                                                                                                                                                                                                         �          �          V       f�S     �         �    �          �      entity somador32 is   
    port (   '        a : in bit_vector(31 downto 0);   '        b : in bit_vector(31 downto 0);   '        r : out bit_vector(31 downto 0)       );   end entity somador32;       'architecture behavioral of somador32 is   +    signal carry : bit_vector(31 downto 0);   begin   "    sum: for i in 0 to 30 generate   +        r(i) <= A(i) xor B(i) xor carry(i);   T        carry(i+1) <= (A(i) and B(i)) or (A(i) and carry(i)) or (B(i) and carry(i));       end generate;       +    r(31) <= A(31) xor B(31) xor carry(31);          end architecture behavioral;    5��                                                 5�_�  �          �  �   <       ����                                                                                                                                                                                                                                                                                                                �          =   .       =   /       V   9    f�(     �   ;   =         5��    ;           Y           �      Y               5�_�  �  �      �  �   6        ����                                                                                                                                                                                                                                                                                                                E           �          �   %       V   9    f<@     �   5   7        5��    5                      W                     5�_�  �  �          �   5        ����                                                                                                                                                                                                                                                                                                                D           �          �   %       V   9    f<B     �   4   6        5��    4                      I                     5�_�  �              �   5        ����                                                                                                                                                                                                                                                                                                                C           �          �   %       V   9    f<B   E �   4   6        5��    4                      I                     5�_�  �  �      �  �  %   !    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6L     �  $  &  5      ,            elsif (iteration = 63) and  then5��    $  !                  @!                     �    $  %                  D!                     �    $  $                 C!                    5�_�  �  �          �  %   '    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6Q     �  $  &  5      .            elsif (iteration = 63) and () then5��    $  '                  F!                     5�_�  �              �  %   (    ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f6Q     �  $  &  5      6            elsif (iteration = 63) and (done = 0) then5��    $  (                  G!                     �    $  *                 I!                    �    $  .                 M!                    5�_�  �          �  �  '       ����                                                                                                                                                                                                                                                                                                                F           �   ,          ,          ,    f5�     �  '  (  .    �  &  ,  .      +                haso <= haso(31 downto 0));   +            end if;     haso(63 downto 32))   +        end if;         haso(95 downto 64))   +                        haso(127 downto 96)       end process;5��    &                    z!                     �    '                    �!                     �    (                    �!                     �    )                  +   �!              +       5��