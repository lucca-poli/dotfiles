Vim�UnDo� �2��p�=�j}�lq��h��bs�!��M   3   .        d2 : out std_logic_vector(3 downto 0);   
   	                       fs     _�                            ����                                                                                                                                                                                                                                                                                                                                                             fst     �                $architecture arch of contador_bcd is�         3      entity contador_bcd is 5��                        M                     �                        �                    5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                             fs�     �   	      3      6        primeiro_d : out std_logic_vector(3 downto 0);5��    	          
          �       
              5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             fs�     �   
      3      5        segundo_d : out std_logic_vector(3 downto 0);5��    
          	                	              5�_�      
                     ����                                                                                                                                                                                                                                                                                                                                                             fs�     �         3      6        terceiro_d : out std_logic_vector(3 downto 0);5��              
          4      
              5�_�                
   0       ����                                                                                                                                                                                                                                                                                                                                                             fs�     �   /   1   3      +    digito2 <= std_logic_vector(signal_d2);5��    /                    �                    5�_�   
                 1       ����                                                                                                                                                                                                                                                                                                                                                             fs�     �   0   2   3      +    digito1 <= std_logic_vector(signal_d1);5��    0                                         5�_�                    2       ����                                                                                                                                                                                                                                                                                                                                                             fs�     �   1   3   3      +    digito0 <= std_logic_vector(signal_d3);5��    1                    G                    5�_�                    2       ����                                                                                                                                                                                                                                                                                                                                                             fs�    �   1   3   3      &    d0 <= std_logic_vector(signal_d3);5��    1                    H                    5�_�                   
   	    ����                                                                                                                                                                                                                                                                                                                            
   	          	          	    fs     �   	      3      .        d1 : out std_logic_vector(3 downto 0);   .        d2 : out std_logic_vector(3 downto 0);   .        d3 : out std_logic_vector(3 downto 0);5��    	   	                 �                     �    
   	                                     �       	                 5                    5�_�                     0       ����                                                                                                                                                                                                                                                                                                                            0          2                 fs    �   /   3   3      &    d3 <= std_logic_vector(signal_d2);   &    d2 <= std_logic_vector(signal_d1);   &    d1 <= std_logic_vector(signal_d3);5��    /                    �                    �    0                    !                    �    1                    H                    5�_�                   
   	    ����                                                                                                                                                                                                                                                                                                                            
   	          	          	    fs     �   	      3      .        d2 : out std_logic_vector(3 downto 0);   .        d3 : out std_logic_vector(3 downto 0);   .        d4 : out std_logic_vector(3 downto 0);5��    	   	                 �                     �    
   	                                     �       	                 5                    5�_�                     
   	    ����                                                                                                                                                                                                                                                                                                                            
   	          	          	    fs     �   	      3      -        d : out std_logic_vector(3 downto 0);5��    	   	                  �                      5�_�             
      0       ����                                                                                                                                                                                                                                                                                                                                                             fs�     �   /   1   3      &    d2 <= std_logic_vector(signal_d2);5��    /                    �                    5�_�      	              1       ����                                                                                                                                                                                                                                                                                                                                                             fs�     �   0   2   3      &    d1 <= std_logic_vector(signal_d1);5��    0                                         5�_�                 	   2       ����                                                                                                                                                                                                                                                                                                                                                             fs�     �   1   3   3      &    d0 <= std_logic_vector(signal_d3);5��    1                    G                    5�_�              	      2       ����                                                                                                                                                                                                                                                                                                                                                             fs�     �   1   3   3      &    d0 <= std_logic_vector(signal_d3);5��    1                    G                    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             fs[     �         3      entity contador_3dig is 5��                        V                     5��