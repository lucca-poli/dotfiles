Vim�UnDo� �I-/�]O�	�Ɇ���P"������.}�   `   1    q <= (x ror 2) xor (x ror 13) xor (x ror 22);   "                         e�P�    _�                        	    ����                                                                                                                                                                                                                                                                                                                                                             e�OE    �         _      use IEEE.NUMERIC_BIT.ALL;5��       	                                      �       	                                      �       	                                      �       	                                      5�_�                           ����                                                                                                                                                                                                                                                                                                                            B           >           V        e�P�     �         `       �         _    5��                          (                      �                          (                      �                         -                      �                        ,                     �                         -                      �                        ,                     �                         -                      �                        ,                     �                         -                      �                        ,                     �                        ,                     �                        ,                     �              
           -       
               �                        ,                     �                        ;                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            C           ?           V        e�P�    �         `      use.numeric_std.all;5��                        +                     5�_�                     "       ����                                                                                                                                                                                                                                                                                                                            C           ?           V        e�P�     �   !   #   `      3    q <= (x ror 2) s xor (x ror 13) xor (x ror 22);5��    !                                          �    !                                          �    !                                          5��