Vim�UnDo� 1�m�{>Z{'X�<�+E����m�.nι[���   0   entity contador_m is                             fs�    _�                             ����                                                                                                                                                                                                                                                                                                                                                  V        fs�    �                 B------------------------------------------------------------------   -- Arquivo   : contador_m.vhd   <-- Projeto   : Experiencia 2 - Comunicacao Serial Assincrona   B------------------------------------------------------------------   !-- Descricao : contador binario     0--             > parametro M: modulo de contagem   5--             > parametro N: numero de bits da saida   --   8--             saidas fim de contagem e meio de contagem   --   B------------------------------------------------------------------   -- Revisoes  :   6--     Data        Versao  Autor             Descricao   ;--     09/09/2021  1.0     Edson Midorikawa  versao inicial   >--     31/08/2022  2.0     Edson Midorikawa  revisao do codigo   4--     04/09/2022  2.1     Edson Midorikawa  revisao   B------------------------------------------------------------------    5��                                   &              5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        fs�    �                -architecture contador_m_arch of contador_m is�                end entity contador_m;�         0      entity contador_m is5��              
          M       
              �              
          �      
              �              
          �      
              �       '       
          �      
              5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        fs�     �         0      entity contador_ is5��                         V                      5��