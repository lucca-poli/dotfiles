Vim�UnDo� ��B�����șo�$'�A�d��L���xR�U                                      e�G�    _�                             ����                                                                                                                                                                                                                                                                                                                                                             e�F�     �                   5��                                                  �                                                �                                                �                                                �                                                5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             e�F�     �                  dawd5��                                                  5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             e�F�     �                   5�5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             e�F�     �                   5��                                                  5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�F�     �                  �               5��                                                �                                                �                                                �                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�G      �                dawdlj5��                                                5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             e�G     �                  5��                                                  5�_�      	                      ����                                                                                                                                                                                                                                                                                                                                                             e�G     �                 5��                                                5�_�      
           	           ����                                                                                                                                                                                                                                                                                                                                                             e�G     �                 kdwjadkjwakd    5��                                                5�_�   	              
           ����                                                                                                                                                                                                                                                                                                                                                             e�G_     �                 use IEEE.numeric_std.all;�                   5��                                                  �        
                  
                      �        	                  	                      �                                              �                                              �                                              �                                                �                                        D       �                          L                       5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                             e�Gf     �                use IEEE.std_logic_1164.all;   use IEEE.numeric_std.all;5��                                 7               5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             e�Gh     �                 use IEEE.numeric_std.all;�                  library library IEEE;5��                                                �                                                �                                                �                                                �                                                �                                                �                                                  �                                          D       �                         D                      �                         D                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             e�G     �                use IEEE.std_logic_1164.all;   use IEEE.numeric_std.all;5��                                 7               5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             e�G�    �                 library IEEE;5��                                                5��