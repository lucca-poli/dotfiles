Vim�UnDo�  ��|��V���}}���|@�T	Z���S�}]   �       signal    g         �       �   �   �    fC��    _�                           ����                                                                                                                                                                                                                                                                                                                            n          q           V       f;Q�     �         �              �         �    5��                          e               	       �                         m                      �                         r                      �                         q                      �                         p                      �       
                  o                      �       	                  n                      �                     	   m              	       �              	          m       	              �                     
   m              
       �                        v                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            o          r           V       f;Q�     �         �              WIDTH: natural := 75��                         d                      �                        d                     5�_�                           ����                                                                                                                                                                                                                                                                                                                            o          r           V       f;Q�     �         �              STOP_BITS := 25��                         w                      �                        {                     5�_�      "              B       ����                                                                                                                                                                                                                                                                                                                            o          r           V       f;Q�    �   A   B          %    constant STOP_BITS: natural := 3;5��    A                      ]      &               5�_�      #           "   8        ����                                                                                                                                                                                                                                                                                                                            n          q           V       f;S�     �   s   u          -                            state <= sending;�   q   s          #                    when sending =>�   n   p          )                        state <= sending;�   7   9   �      ;    type transmiter is (starting, sending, stopping, idle);5��    7   "              	                	       �    n   !              	   ]             	       �    q                 	   �             	       �    s   %              	                	       5�_�   "   $           #   ?        ����                                                                                                                                                                                                                                                                                                                            n          q           V       f;S�     �   �   �          \                        if stop_bits_sent < STOP_BITS then -- numero de stop bits arbitrario�   t   v          >                            if signal_bits_sent = WIDTH-1 then�   r   t          8                        if signal_bits_sent < WIDTH then�   O   Q          H        port map(new_clk, reset, start_stop, done_stop, stop_bits_sent);�   K   M          N        port map(new_clk, reset, start_signal, done_signal, signal_bits_sent);�   >   @   �      5    signal signal_bits_sent, stop_bits_sent: natural;5��    >                    #                    �    >   +                 7                    �    K   H                 ^                    �    O   B                                     �    r   '                 �                    �    t   +                 d                    �    �   %                 b                    5�_�   #   %           $   g   %    ����                                                                                                                                                                                                                                                                                                                            n          q           V       f;S�     �   f   h   �      .                            state <= starting;5��    f   %                 t
                    �    f   +                  z
                     �    f   *                  y
                     �    f   )                  x
                     �    f   (                  w
                     �    f   '                  v
                     �    f   &                  u
                     �    f   %                 t
                    �    f   (                  w
                     �    f   '                  v
                     �    f   &                  u
                     �    f   %              	   t
             	       �    f   %       	          t
      	              �    f   %              	   t
             	       5�_�   $   &           %   p   +    ����                                                                                                                                                                                                                                                                                                                            n          q           V       f;T     �   o   p          ,                        start_signal <= '0';5��    o                      y      -               5�_�   %   '           &   q        ����                                                                                                                                                                                                                                                                                                                            n          p           V       f;T     �   q   s   �    �   q   r   �    5��    q                      �              -       5�_�   &   (           '   n       ����                                                                                                                                                                                                                                                                                                                            n          p           V       f;T     �   m   n          $                    when starting =>   +                        state <= receiving;5��    m                      (      Q               5�_�   '   )           (   n        ����                                                                                                                                                                                                                                                                                                                            n          n           V       f;T     �   m   n           5��    m                      (                     5�_�   (   *           )   K       ����                                                                                                                                                                                                                                                                                                                            n          n           V       f;T<     �   J   L   �              generic map(WIDTH+1)5��    J                                          �    J                                          5�_�   )   +           *   �       ����                                                                                                                                                                                                                                                                                                                            n          n           V       f;U,     �   �   �   �      (                            done <= '1';5��    �                     �                     5�_�   *   ,           +   �       ����                                                                                                                                                                                                                                                                                                                            n          n           V       f;U-     �   �   �   �      *                            state <= idle;5��    �                                          5�_�   +   -           ,   �       ����                                                                                                                                                                                                                                                                                                                            n          n           V       f;U1     �   �   �   �                                  �   �   �   �    5��    �                      �              !       �    �                   #   �              #       �    �   "                  �                     �    �   !                  �                     �    �                      �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�   ,   .           -   �   -    ����                                                                                                                                                                                                                                                                                                                            n          n           V       f;U8     �   �   �   �      -                            if serial_data = 5��    �   -                  �                     5�_�   -   /           .   �   .    ����                                                                                                                                                                                                                                                                                                                            n          n           V       f;U9     �   �   �   �      /                            if serial_data = ''5��    �   .                  �                     5�_�   .   0           /   �   0    ����                                                                                                                                                                                                                                                                                                                            n          n           V       f;U;     �   �   �   �      0                            if serial_data = '1'5��    �   0                  �                     5�_�   /   1           0   �   1    ����                                                                                                                                                                                                                                                                                                                            n          n           V       f;U?     �   �   �   �      %                                state�   �   �   �                                       �   �   �   �    5��    �                                    !       �    �                      ?                     �    �   "                  A                     �    �   !                 @                    �    �                                           �    �                     ?                     �    �                  #   @             #       �    �   "                  b                     �    �   !                  a                     �    �                  
   `             
       �    �   )                  i                     �    �   (                  h                     �    �   '                  g                     �    �   &                  f                     �    �   %                  e                     �    �   $                  d                     �    �   #                  c                     �    �   "                  b                     �    �   !                  a                     �    �                     `                    �    �   $                  d                     �    �   #                  c                     �    �   "                  b                     �    �   !                  a                     �    �                     `                    �    �                     `                    �    �                     `                    �    �   ,                  l                     �    �   +                  k                     �    �   *                  j                     �    �   )                 i                    �    �   ,                  l                     �    �   +                  k                     �    �   *                  j                     �    �   )              	   i             	       �    �   )       	          i      	              �    �   )              
   i             
       5�_�   0   2           1   �        ����                                                                                                                                                                                                                                                                                                                            i   %       k   .       V   2    f;UX     �   �   �   �    5��    �                      t              !       �    �                       t                      5�_�   1   3           2   �        ����                                                                                                                                                                                                                                                                                                                            i   %       k   .       V   2    f;UY     �   �   �   �    �   �   �   �    5��    �                      u              �       5�_�   2   4           3   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f;U[     �   �   �   �      0                            start_signal <= '1';   .                            shift_data <= '1';�   �   �   �      &                            -- Control5��    �                     �                     �    �                     �                     �    �                     �                     5�_�   3   5           4   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f;U^    �   �   �   �                                       �   �   �   �    5��    �                                    !       �    �                      (                     �    �                                           �    �                      (                     5�_�   4   6           5   8       ����                                                                                                                                                                                                                                                                                                                            �          �                 f;Uq     �   7   9   �      =    type transmiter is (starting, receiving, stopping, idle);5��    7                                          5�_�   5   7           6   8       ����                                                                                                                                                                                                                                                                                                                            �          �                 f;Ur    �   7   9   �      5    type transmiter is (, receiving, stopping, idle);5��    7                                          5�_�   6   ;           7   p   7    ����                                                                                                                                                                                                                                                                                                                            �          �                 f;Vt     �   o   q   �      <                        if signal_bits_received < WIDTH then5��    o   7                  �                     5�_�   7   <   8       ;   r   <    ����                                                                                                                                                                                                                                                                                                                            �          �                 f;V�    �   q   s   �      B                            if signal_bits_received = WIDTH-1 then5��    q   <                                     5�_�   ;   =           <   �        ����                                                                                                                                                                                                                                                                                                                            �          �   #       V   <    f;We     �   �   �                                       else   3                                state <= receiving;       *                                -- Control   4                                start_signal <= '1';   2                                shift_data <= '1';   #                            end if;5��    �                                          5�_�   <   >           =   �       ����                                                                                                                                                                                                                                                                                                                            �          �   #       V   <    f;Wh     �   �   �          5                            if serial_data = '1' then5��    �                      �      6               5�_�   =   ?           >   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   f;Wm     �   �   �   �      ,                                done <= '1';5��    �                     �                     5�_�   >   @           ?   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   f;Wo     �   �   �   �      .                                state <= idle;5��    �                                          5�_�   ?   A           @   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   f;Wq     �   �   �   �      *                                -- Control5��    �                     /                     5�_�   @   B           A   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   f;Wr     �   �   �   �      4                                start_signal <= '0';5��    �                     V                     5�_�   A   C           B   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   f;Wr     �   �   �   �      2                                start_stop <= '0';5��    �                     �                     5�_�   B   D           C   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   f;Ws     �   �   �   �      2                                shift_data <= '0';5��    �                     �                     5�_�   C   E           D   k       ����                                                                                                                                                                                                                                                                                                                            �           �                   f;X�     �   j   k          .                            shift_data <= '1';5��    j                      �
      /               5�_�   D   F           E   p       ����                                                                                                                                                                                                                                                                                                                            �           �                   f;X�     �   p   r   �    �   p   q   �    5��    p                      �              /       5�_�   E   G           F   r   5    ����                                                                                                                                                                                                                                                                                                                            �           �                   f;Yj     �   q   s   �      B                            if signal_bits_received = WIDTH-2 then5��    q   4                                     5�_�   F   H           G   r   <    ����                                                                                                                                                                                                                                                                                                                            �           �                   f;Y�     �   q   s   �      B                            if signal_bits_received < WIDTH-2 then5��    q   <                                     5�_�   G   I           H   r   <    ����                                                                                                                                                                                                                                                                                                                            �           �                   f;Y�     �   q   r          B                            if signal_bits_received < WIDTH-1 then5��    q                      �      C               5�_�   H   J           I   s   "    ����                                                                                                                                                                                                                                                                                                                            �           �                   f;Y�     �   r   s          #                            end if;5��    r                            $               5�_�   I   K           J   r        ����                                                                                                                                                                                                                                                                                                                            �           �                   f;Y�     �   q   s   �      2                                shift_data <= '0';5��    q                     �                     5�_�   J   L           K   r       ����                                                                                                                                                                                                                                                                                                                            �           �                   f;Y�     �   q   r          .                            shift_data <= '0';5��    q                      �      /               5�_�   K   N           L   t       ����                                                                                                                                                                                                                                                                                                                                       �                   f;Y�    �   t   v   �    �   t   u   �    5��    t                      Y              /       5�_�   L   O   M       N   v        ����                                                                                                                                                                                                                                                                                                                            v           x           V        f;ZZ     �   u   v          #                            -- Data   Q                            parity_bit <= not data_to_parity(word); -- parity bit   2                            parallel_data <= word;5��    u                      �      �               5�_�   N   P           O   {        ����                                                                                                                                                                                                                                                                                                                            v           v           V        f;Z_     �   {   }   �    5��    {                      �                     �    {                      �                     5�_�   O   Q           P   |        ����                                                                                                                                                                                                                                                                                                                            v           v           V        f;Z_    �   |   �   �    �   |   }   �    5��    |                      �              �       5�_�   P   R           Q   q       ����                                                                                                                                                                                                                                                                                                                            v           v           V        f;]L     �   p   q          .                            shift_data <= '1';5��    p                      �      /               5�_�   Q   S           R   j       ����                                                                                                                                                                                                                                                                                                                            u           u           V        f;]R   	 �   j   l   �    �   j   k   �    5��    j                      �
              /       5�_�   R   T           S      *    ����                                                                                                                                                                                                                                                                                                                            �          �           v        fC��     �      �   �                                  �      �   �    5��                          7                     �                         S                     �       !                  X                     �                          W                     �                        V                    �       $                  [                     �       #                  Z                     �       "                  Y                     �       !                  X                     �                          W                     �                        V                    �                        V                    �                        V                    �       7                  n                     �       6                  m                     �       5                  l                     �       4              	   k             	       �       4       	          k      	              �       4                 k                    �       @                 w                    �       @                 w                    �       @                 w                    �       D                 {                     �    �                  (   |             (       5�_�   S   U           T   �   (    ����                                                                                                                                                                                                                                                                                                                            �          �           v        fC��     �   �   �   �      (                                done <= 5��    �   (                  �                     5�_�   T   V           U   �   *    ����                                                                                                                                                                                                                                                                                                                            �          �           v        fC�      �   �   �   �      *                                done <= ''5��    �   )                 �                    5�_�   U   W           V   �   %    ����                                                                                                                                                                                                                                                                                                                            �          �           v        fC�     �   �   �   �      (                            done <= '1';5��    �   %                 �                    5�_�   V   X           W   �       ����                                                                                                                                                                                                                                                                                                                            �          �           v        fC�	   
 �   �   �   �                                       �   �   �   �    5��    �                      �                     �    �                  $   �             $       �    �                      �                     �    �                      �                     5�_�   W   Y           X   B       ����                                                                                                                                                                                                                                                                                                                            �          �           v        fC�9     �   A   C   �          signal new_clk: bit;5��    A                 
   h             
       5�_�   X   d           Y   H        ����                                                                                                                                                                                                                                                                                                                            H          Z          V       fC�O     �   V   X          $        if rising_edge(new_clk) then�   T   V              process(new_clk) is�   R   T          @        port map(reset, new_clk, shift_data, serial_data, word);�   O   Q          L        port map(new_clk, reset, start_stop, done_stop, stop_bits_received);�   K   M          R        port map(new_clk, reset, start_signal, done_signal, signal_bits_received);�   G   I   �      !        port map(clock, new_clk);5��    G                    �                    �    K                    !                    �    O                    �                    �    R                    G                    �    T                    �                    �    V                    �                    5�_�   Y   e   Z       d   �       ����                                                                                                                                                                                                                                                                                                                            H          Z          V       fC��     �   �   �          (                            done <= '0';5��    �                      �      )               5�_�   d   f           e   F       ����                                                                                                                                                                                                                                                                                                                            F          F          v       fC��     �   E   G   �          clocking: slow_clk5��    E                    �                    5�_�   e   g           f          ����                                                                                                                                                                                                                                                                                                                            F          F          v       fC��     �          �    5��                                                  5�_�   f   h           g           ����                                                                                                                                                                                                                                                                                                                            G          G          v       fC��     �       	   �    �         �    5��                                           �       5�_�   g   i           h      !    ����                                                                                                                                                                                                                                                                                                                            O          O          v       fC��     �         �      !        rst, clk, enable: in bit;5��       !                 g               	       �                         h                     5�_�   h   j           i          ����                                                                                                                                                                                                                                                                                                                            P          P          v       fC��     �         �              sample: out bit;5��                                               5�_�   i   k           j   	       ����                                                                                                                                                                                                                                                                                                                            P          P          v       fC�     �         �      end architecture �   
      �      architecture rtl of  is�         �          �   
      �      arch�   	      �       �   	      �    5��    	                      �                      �    	                      �                      �    
                      �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                     �    
                     �                     �    
                     �                     �    
                     �                     �    
                    �                      �                          �                       �                        �                      �                         �                      �    
                     �                      �                         �                      5�_�   j   l           k          ����                                                                                                                                                                                                                                                                                                                                                v       fC�     �         �    �         �      end architecture rtl;�   
      �      )architecture Behavioral of tx_receptor is�         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �         �    �   
      �      "architecture rtl of tx_receptor is5��    
                    �                     �                        �                     �    
                     �                      �                        �                     �    
                     �                      �                        �                     �    
                     �                      �                        �                     �    
                     �                      �                        �                     �    
                     �                      �                        �                     �    
                     �                      �                        �                     �    
                     �                      �                        �                     �    
                     �                      �                        �                     �    
                     �                      �                        �                     �    
                     �                      �                        �                     �    
                     �                      �                        �                     �    
                     �                      �    
                 
   �              
       �    
          
          �       
              �    
                 
   �              
       �                     
   �              
       5�_�   k   m           l          ����                                                                                                                                                                                                                                                                                                                               %                 v       fC�
     �   
      �      )architecture Behavioral of tx_receptor is5��    
                    �                     �    
                      �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                     �                      �    
                    �                     �    
                    �                     �    
                    �                     5�_�   l   n           m          ����                                                                                                                                                                                                                                                                                                                               %                 v       fC�-     �         �          �         �    5��                          �                      �                          �                      �                         �                      �                         �                      �                         �                      �                         �                      �                         �                      �                        �                     5�_�   m   o           n          ����                                                                                                                                                                                                                                                                                                                            i           �           V        fC�v     �      K   �    �         �    5��                   :       �               �      5�_�   n   p           o          ����                                                                                                                                                                                                                                                                                                                            �           �           V        fC�     �         �          process(slowed_clk) is5��              
                 
              5�_�   o   q           p          ����                                                                                                                                                                                                                                                                                                                            �           �           V        fC��     �         �      '        if rising_edge(slowed_clk) then5��              
          )      
              5�_�   p   r           q           ����                                                                                                                                                                                                                                                                                                                                                V       fC��     �         �      )                state <= idle; -- repouso�                                done <= '0';                       -- Control   $                start_signal <= '0';   "                start_stop <= '0';   "                shift_data <= '0';5��                          }      �               �                        c                    �                         e                     �                         d                     �                        c                    �                        c                    �                        c                    5�_�   q   s           r          ����                                                                                                                                                                                                                                                                                                                                                V       fC��     �         �                  if reset = '1' then5��                        B                    5�_�   r   t           s           ����                                                                                                                                                                                                                                                                                                                                      B          V       fC��    �         �                          offset�         �                      case state is�             +                            when idle =>   $                        done <= '0';       1                        if serial_data = '0' then   /                            state <= receiving;       &                            -- Control   0                            start_signal <= '1';   .                            shift_data <= '1';                           end if;       %                    when receiving =>   ,                        start_signal <= '0';   >                        if signal_bits_received < WIDTH-1 then   /                            state <= receiving;                           else   .                            state <= stopping;   .                            start_stop <= '1';   .                            shift_data <= '0';                           end if;       $                    when stopping =>   `                        if stop_bits_received < STOP_BITS then -- numero de stop bits arbitrario   .                            state <= stopping;   .                            start_stop <= '0';       #                            -- Data   Q                            parity_bit <= not data_to_parity(word); -- parity bit   2                            parallel_data <= word;   D                            if stop_bits_received = STOP_BITS-1 then   ,                                done <= '1';   #                            end if;                           else   *                            state <= idle;       &                            -- Control   0                            start_signal <= '0';   .                            start_stop <= '0';   .                            shift_data <= '0';                           end if;                   end case;               end if;5��           +               �      Q              �                        �                    �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    �                        �                    �                        �                    �                        �                    �       "                 �                     �                         �                    �                         �                     �                        �                    �                        �                    �                        �                    �                         �                     �                         �                     5�_�   s   u           t          ����                                                                                                                                                                                                                                                                                                                                                V       fC��     �         �                          offse5��                         �                     �                          �                     �                         �                     �                        �                    �                        �                    �                     	   �             	       �       &                 �                    �       )                 �                     �                        �                    �                         �                     �                        �                     �                         �                    �                          �                     5�_�   t   v           u          ����                                                                                                                                                                                                                                                                                                                                                V       fC�,     �         �                      offset <= 3;5��                        k                    5�_�   u   w           v      %    ����                                                                                                                                                                                                                                                                                                                                                V       fC�7     �         �      )                    offset <= offset - 1;5��       %                 �                    5�_�   v   x           w          ����                                                                                                                                                                                                                                                                                                                                                V       fC�I     �         �      "                if offset > 0 then5��                        �                    5�_�   w   y           x          ����                                                                                                                                                                                                                                                                                                                                                V       fC�]     �         �      "                if offset < 0 then5��                        �                    5�_�   x   {           y          ����                                                                                                                                                                                                                                                                                                                                                V       fC�w     �         �           signal offset: natural := 3;5��                        �                     5�_�   y   |   z       {           ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �                )                    offset <= offset + 1;�                "                if offset < 4 then�                                offset <= 0;�         �           signal offset: natural := 0;5��                        �                     �                        b                    �                        �                    �                        �                    �                        �                    5�_�   {   }           |          ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �                              sample�         �                          �         �    5��                          �                     �                         �                     �       #                 �                    �       #                 �                    �       #                 �                    �       '                 �                     �                         �                    �                                              �                                              �                                              �                                              �                                            �                                            �                                            �                                            5�_�   |   ~           }      "    ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �      "                        sample <= 5��       "                                       5�_�   }              ~      #    ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �      $                        sample <= ''5��       #                                       5�_�   ~   �                 %    ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �      %                        sample <= '1'5��       %                                       5�_�      �           �           ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �       5��                          5                     �                         L                     �                         K                     �                         J                     �                        I                    �                        I                    �                        I                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �                          counter <= 5��                         T                     5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �      !                    counter <= ''5��                          U                     5�_�   �   �           �      "    ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �      "                    counter <= '0'5��       "                  W                     5�_�   �   �           �      "    ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �    �         �    5��                          Y              $       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �      #                    counter <= '0';5��                        m                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �                          �         �    5��                          |                     �                         �                     �                         |                    �                         �                     �                         �                     �                        �                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �                              �         �    5��                                                �                         8                     �                                              �                         8                     �                        :                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �      !   �                      �      !   �    5��                          �                     �                         �                     �                         �                    �                         �                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �      #                    counter <= '0';5��                         p                     5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �      "                    counter <= 0';5��                          q                     5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �         �      !        rst, clk, enable: in bit;5��                         X                      5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                  V        fC��    �         �              rst, clk, : in bit;5��                         V                      5�_�   �   �           �   l       ����                                                                                                                                                                                                                                                                                                                                                  V        fC�	     �   k   m   �          clocking: sample_clk5��    k          
          �	      
              5�_�   �   �           �   m       ����                                                                                                                                                                                                                                                                                                                                                  V        fC�     �   l   m          		generic map(1)5��    l                      �	                     5�_�   �   �           �   m       ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �   l   n   �      $        port map(clock, slowed_clk);5��    l                     �	                     5�_�   �   �           �   h        ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �   {   }          '        if rising_edge(slowed_clk) then�   y   {              process(slowed_clk) is�   w   y          C        port map(reset, slowed_clk, shift_data, serial_data, word);�   t   v          O        port map(slowed_clk, reset, start_stop, done_stop, stop_bits_received);�   p   r          U        port map(slowed_clk, reset, start_signal, done_signal, signal_bits_received);�   l   n          &        port map(, clock, slowed_clk);�   g   i   �          signal slowed_clk: bit;5��    g                    k	                    �    l                    �	                    �    p                    
                    �    t                    �
                    �    w                    :                    �    y                    s                    �    {                    �                    5�_�   �   �           �   f       ����                                                                                                                                                                                                                                                                                                                                                  V        fC�R     �   f   h   �          �   f   h   �    5��    f                      _	                     �    f                     c	                     5�_�   �   �           �   {       ����                                                                                                                                                                                                                                                                                                                                                  V        fC�Y     �   z   |   �          process(sample_clk) is5��    z          
                
              5�_�   �   �           �   }       ����                                                                                                                                                                                                                                                                                                                                                  V        fC�\     �   |   ~   �      '        if rising_edge(sample_clk) then5��    |          
          �      
              5�_�   �   �           �   n       ����                                                                                                                                                                                                                                                                                                                                                  V        fC��     �   m   o   �      &        port map(, clock, sample_clk);5��    m                     �	                     �    m                    �	                    �    m                    �	                    5�_�   �               �   g       ����                                                                                                                                                                                                                                                                                                                                                  V        fC��    �   f   h   �          signal 5��    f                     j	                     �    f                    k	                    �    f                     l	                     �    f                     k	                     �    f                    j	                    �    f                    j	                    �    f                    j	                    5�_�   y           {   z           ����                                                                                                                                                                                                                                                                                                                                                V       fC�~     �              �         �       5��                          �       �               �                           �                       5�_�   Y   [       d   Z   �       ����                                                                                                                                                                                                                                                                                                                            H          Z          V       fC��     �   �   �        5��    �                      �      -               5�_�   Z   \           [   u       ����                                                                                                                                                                                                                                                                                                                            H          Z          V       fC��     �   u   v   �    �   u   v   �      ,                                done <= '1';5��    u                      �              -       5�_�   [   ]           \   v        ����                                                                                                                                                                                                                                                                                                                            H          Z          V       fC��     �   u   w   �      (                            done <= '1';5��    u                     �                     5�_�   \   ^           ]   y       ����                                                                                                                                                                                                                                                                                                                            H          Z          V       fC��     �   y   z   �                              �   y   {   �                              donw               d5��    y                                           �    y                                         �    y                    (                     �    z                    9                    �    z                    5                    5�_�   ]   _           ^   {       ����                                                                                                                                                                                                                                                                                                                            H          Z          V       fC�     �   z   |        5��    z                      )                     5�_�   ^   `           _   z       ����                                                                                                                                                                                                                                                                                                                            H          Z          V       fC�     �   y   {   �                               done <= 5��    y                    '                    5�_�   _   a           `   z        ����                                                                                                                                                                                                                                                                                                                            H          Z          V       fC�     �   y   {   �      "                        done <= ''5��    y                      ,                     5�_�   `   b           a   z   !    ����                                                                                                                                                                                                                                                                                                                            H          Z          V       fC�     �   y   {   �      #                        done <= '0'5��    y   !                  -                     5�_�   a   c           b   z   #    ����                                                                                                                                                                                                                                                                                                                            H          Z          V       fC�     �   y   {   �      $                        done <= '0';5��    y   #                  /                     5�_�   b               c   z   #    ����                                                                                                                                                                                                                                                                                                                            H          Z          V       fC�!     �   y   {        5��    y                            %               5�_�   L           N   M   v        ����                                                                                                                                                                                                                                                                                                                            v          v          V       f;ZF     �   u   y        5��    u                      �      �               5�_�   7   9       ;   8   r   8    ����                                                                                                                                                                                                                                                                                                                            �          �                 f;Vz     �   q   s        5��    q                      �      C               5�_�   8   :           9   s   "    ����                                                                                                                                                                                                                                                                                                                            �          �                 f;V|     �   r   t        5��    r                            $               5�_�   9               :   r        ����                                                                                                                                                                                                                                                                                                                            �          �                 f;V}     �   q   s   �      .                            shift_data <= '0';5��    q                     �                     5�_�      !       "       g   %    ����                                                                                                                                                                                                                                                                                                                            n          q           V       f;S�     �   f   h   �      &                            state <= ;5��    f   %                  b
                     5�_�                   !   g   %    ����                                                                                                                                                                                                                                                                                                                            n          q           V       f;S�     �   f   h   �      '                            state <= s;5��    f   %                  b
                     5�_�                    g   %    ����                                                                                                                                                                                                                                                                                                                                                             f:�
     �   f   h   �      -                            state <= sending;5��    f   %                 g
                    5�_�                    p   +    ����                                                                                                                                                                                                                                                                                                                                                             f:�     �   o   q        5��    o                      h      -               5�_�                    r        ����                                                                                                                                                                                                                                                                                                                                                             f:�$     �   r   s   �    �   q   r   �      ,                        start_signal <= '0';5��    q                      �              -       5�_�                    7        ����                                                                                                                                                                                                                                                                                                                                                             f:�E     �   6   8   �      =    type transmiter is (starting, receiving, stopping, idle);�   f   h          /                            state <= receiving;�   n   p          +                        state <= receiving;�   p   r          %                    when receiving =>�   s   u          /                            state <= receiving;5��    6   "              	   �             	       �    f   %              	   i
             	       �    n   !              	   c             	       �    p                 	   �             	       �    s   %              	                 	       5�_�                   >        ����                                                                                                                                                                                                                                                                                                                                                             f:�|     �   =   ?   �      =    signal signal_bits_received, stop_bits_received: natural;�   K   M          R        port map(new_clk, reset, start_signal, done_signal, signal_bits_received);�   O   Q          L        port map(new_clk, reset, start_stop, done_stop, stop_bits_received);�   r   t          <                        if signal_bits_received < WIDTH then�   t   v          B                            if signal_bits_received = WIDTH-1 then�   �   �          `                        if stop_bits_received < STOP_BITS then -- numero de stop bits arbitrario5��    =                                        �    =   +                                     �    K   H                 c                    �    O   B                 
                    �    r   '                 �                    �    t   +                 j                    �    �   %                 h                    5�_�                    n        ����                                                                                                                                                                                                                                                                                                                            n          n           V       f:��     �   m   q        5��    m                      -      R               5�_�      	              7       ����                                                                                                                                                                                                                                                                                                                            n          n           V       f:��     �   6   8   �      5    type transmiter is (, receiving, stopping, idle);5��    6                     �                     5�_�      
           	   7       ����                                                                                                                                                                                                                                                                                                                            n          n           V       f:��     �   6   8   �      3    type transmiter is (receiving, stopping, idle);5��    6                     �                     5�_�   	              
   n       ����                                                                                                                                                                                                                                                                                                                            n          n           V       f:��     �   n   o   �                              �   n   p   �                               done <= 5��    n                      I                     �    n                      I                     5�_�   
                 o        ����                                                                                                                                                                                                                                                                                                                            n          n           V       f:��     �   n   p   �      "                        done <= ''5��    n                      i                     5�_�                    o   !    ����                                                                                                                                                                                                                                                                                                                            n          n           V       f:��     �   n   p   �      #                        done <= '0'5��    n   !                  j                     5�_�                    o   #    ����                                                                                                                                                                                                                                                                                                                            n          n           V       f:��     �   n   p   �      $                        done <= '0';5��    n   #                  l                     5�_�                    �   #    ����                                                                                                                                                                                                                                                                                                                            n          n           V       f:��     �   �   �   �                                  �   �   �   �      -                            if serial_data = 5��    �                      �                     �    �                                          �    �   "                  
                     �    �   !                  	                     �    �                                           �    �                                        �    �                                        �    �                                        5�_�                    �   -    ����                                                                                                                                                                                                                                                                                                                            n          n           V       f:��     �   �   �   �      /                            if serial_data = ''5��    �   -                                       5�_�                    �   .    ����                                                                                                                                                                                                                                                                                                                            n          n           V       f:��     �   �   �   �      0                            if serial_data = '1'5��    �   .                                       5�_�                    �   0    ����                                                                                                                                                                                                                                                                                                                            �          �                 f:��     �   �   �   �      5                            if serial_data = '1' then5��    �   0                                       5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f:��     �   �   �   �      ,                                done <= '1';�   �   �   �      .                                state <= idle;5��    �                     :                     �    �                     g                     5�_�                    �   2    ����                                                                                                                                                                                                                                                                                                                            �          �                 f:��     �   �   �   �      2                                shift_data <= '0';                                else   #                                dwa5��    �   2                  @              !       �    �                      a                     �    �                      A                     �    �                     a                     �    �                  #   b             #       5�_�                    �   "    ����                                                                                                                                                                                                                                                                                                                            �          �                 f:��     �   �   �   �                                       �   �   �   �      #                            end if;5��    �                      �              !       �    �                      �                     �    �                      �                     �    �                      �                     5�_�                    �   "    ����                                                                                                                                                                                                                                                                                                                            �          �                 f:��     �   �   �        5��    �                            -               5�_�                    �   "    ����                                                                                                                                                                                                                                                                                                                            �          �                 f:��     �   �   �   �    �   �   �   �      ,                                done <= '1';5��    �                      �              -       5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f:��     �   �   �   �      (                            done <= '1';5��    �                                          5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            i   %       k   -       V   -    f:�     �   �   �   �      3                                state <= receiving;5��    �                     ~                    �    �   +                  �                     �    �   *                  �                     �    �   )                 �                    �    �   ,                  �                     �    �   +                  �                     �    �   *                  �                     �    �   )                 �                    �    �   0                  �                     �    �   /                  �                     �    �   .                  �                     �    �   -                  �                     �    �   ,                  �                     �    �   +                  �                     �    �   *                  �                     �    �   )              
   �             
       5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            i   %       k   -       V   -    f:�&     �   �   �   �       5��    �                      �              !       �    �                       �                      5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �          �                 f:�'     �   �   �   �    �   �   �   �      &                            -- Control   0                            start_signal <= '1';   .                            shift_data <= '1';5��    �                      �              �       5�_�                     �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f:�)    �   �   �   �      *                                -- Control�   �   �   �      4                                start_signal <= '1';   2                                shift_data <= '1';5��    �                     �                     �    �                     �                     �    �                                          5�_�                    >        ����                                                                                                                                                                                                                                                                                                                                                             f:�f     �   =   ?   �      9    signal signal_bits_received, stop_bits_sent: natural;�   K   M          R        port map(new_clk, reset, start_signal, done_signal, signal_bits_received);�   O   Q          L        port map(new_clk, reset, start_stop, done_stop, stop_bits_received);�   r   t          <                        if signal_bits_received < WIDTH then�   t   v          B                            if signal_bits_received = WIDTH-1 then�   �   �          `                        if stop_bits_received < STOP_BITS then -- numero de stop bits arbitrario5��    =                                        �    K   H                 _                    �    O   B                                     �    r   '                 �                    �    t   +                 f                    �    �   %                 d                    5��