Vim�UnDo� 4�W��ý ��wव��7�}��ޑ�A ����   �                                   f(l�    _�                             ����                                                                                                                                                                                                                                                                                                                                                             f(=I     �                   �               5��                    &                       �      5�_�                    '        ����                                                                                                                                                                                                                                                                                                                                                             f(=s    �   '            �   '            5��    '               $       �              a      5�_�                    &        ����                                                                                                                                                                                                                                                                                                                                       &           V        f(I�     �   &   (   K    5��    &                      �                     5�_�                    '        ����                                                                                                                                                                                                                                                                                                                                       &           V        f(I�    �   '   :   L    �   '   (   L    5��    '                      �              �      5�_�                    &        ����                                                                                                                                                                                                                                                                                                                                                             f(l�     �   '   J   `       �   (   )   `    �   &   )   _       �   &   (   ^    5��    &                      �                     �    &                      �                     �    '               !       �                    5�_�                     I        ����                                                                                                                                                                                                                                                                                                                                                             f(l�    �   H   I           5��    H                      �                     5��