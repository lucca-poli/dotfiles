Vim�UnDo� �SWFv�'�`���J6�/S\V��́�QH�%     $    -- Divisor de clock para 2400 Hz                             f)C�    _�                             ����                                                                                                                                                                                                                                                                                                                                      "          V       f)C�     �              "   I--ENTIDADES AUXILIARES NECESSARIAS---------------------------------------   $    ---Divisor de clock para 9600 Hz   --    library IEEE;   --    use ieee.numeric_bit.all;   --    entity divisorclock4 is   --      Port (   --          clki : in  bit;   --          rst  : in  bit;   --          clko: out bit   
--      );   --    end divisorclock4;   --       *--    architecture arc of divisorclock4 is   c--      constant CLOCK_DIVIDER : integer := 2604; -- 4x mais rapido que o clock de 2400 Hz (9600Hz)   B--      signal counter : unsigned(11 downto 0) := (others => '0');   (--      signal clk_out_int : bit := '0';   --    begin   --      process(clki, rst)   --      begin   --          if rst = '1' then   +--              counter <= (others => '0');   #--              clk_out_int <= '0';   (--          elsif rising_edge(clki) then   3--              if counter = CLOCK_DIVIDER - 1 then   /--                  counter <= (others => '0');   3--                  clk_out_int <= not clk_out_int;   --              else   +--                  counter <= counter + 1;   --              end if;   --          end if;   --      end process;   --       --      clko <= clk_out_int;   --    end architecture;5��            "                       j              5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       f)C�    �               $    -- Divisor de clock para 2400 Hz5��                                              5��