Vim�UnDo� �K�?w���-�ʵ��/�����B��)2�]|   �               reset => reset,   �                      fC��   . _�                            ����                                                                                                                                                                                                                                                                                                                                                             f:kR     �          �      entity sha256_1b is5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f:kS     �          �      entity sha256is5��                                                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f:kW     �         �      end sha256_1b;5��              	          �       	              �       	                 �                     5�_�                    	   !    ����                                                                                                                                                                                                                                                                                                                                                             f:k]     �      
   �      'architecture Behavioral of sha256_1b is5��       !                  �                      5�_�                    	   !    ����                                                                                                                                                                                                                                                                                                                                                             f:k^     �      
   �      #architecture Behavioral of sha256is5��       !                  �                      5�_�                    _   	    ����                                                                                                                                                                                                                                                                                                                                                             f:v�     �   a   c   �              generic�   `   c   �          receiver�   _   b   �              �   _   a   �    5��    _                      �	              	       �    _                      �	                     �    _                     �	              	       �    `                    �	                    �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                    �	                    �    `                    �	                    �    `                    �	                    �    `                     �	                     �    `                     �	                     �    `                    �	                    �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                 
   �	             
       �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                    �	                    �    `   !                  �	                     �    `                      �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                    �	                    �    `   $                  �	                     �    `   #                  �	                     �    `   "                  �	                     �    `   !                  �	                     �    `                      �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                    �	                    �    `   +                  �	                     �    `   *                  �	                     �    `   )                  �	                     �    `   (                  �	                     �    `   '                  �	                     �    `   &                  �	                     �    `   %                  �	                     �    `   $                  �	                     �    `   #                  �	                     �    `   "                  �	                     �    `   !                  �	                     �    `                      �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                     �	                     �    `                    �	                    �    `                    �	                    �    `                    �	                    �    `   ,                 �	                     �    a                     �	                     �    a                    �	                    �    a                    �	                    �    a                    �	                    5�_�                    b       ����                                                                                                                                                                                                                                                                                                                                                             f:v�     �   a   c   �              generic map5��    a                     �	                     5�_�      	              b       ����                                                                                                                                                                                                                                                                                                                                                             f:v�     �   a   c   �              generic map()5��    a                     �	                     5�_�      
           	   b       ����                                                                                                                                                                                                                                                                                                                                                             f:v�     �   a   d   �              generic map(64)5��    a                    �	              	       �    b                     �	                     5�_�   	              
   c       ����                                                                                                                                                                                                                                                                                                                                                             f:v�     �   b   d   �              port map5��    b                     �	                     5�_�   
                 c       ����                                                                                                                                                                                                                                                                                                                                                             f:w	     �   b   d   �              port map()5��    b                     �	                     �    b                     �	                     5�_�                    c       ����                                                                                                                                                                                                                                                                                                                                                             f:w     �   b   e   �              port map(�   c   e                          )�   b   e   �              port map()5��    b                    �	              	       �    c                     �	                    �    b                    �	              	       �    c                     �	                     �    c                      �	                     5�_�                    e       ����                                                                                                                                                                                                                                                                                                                                                             f:w     �   d   f   �                      )5��    d                     �	                     5�_�                    e   	    ����                                                                                                                                                                                                                                                                                                                                                             f:w     �   d   f   �      	        )5��    d   	                  �	                     5�_�                    d        ����                                                                                                                                                                                                                                                                                                                                                             f:w     �   e   i   �      $            enable => done_receiving�   d   g   �                  rst�   c   f   �       5��    c                      �	                     �    c                    �	                    �    c                    �	                    �    c                    �	                    �    c                    �	                    �    c                    
                    �    c                    
                    �    c                    
                    �    c                    
                    �    c                    
                    �    c                    
                    �    c                    
                    �    c                    
                    �    c                    
                    �    c                     
                     �    d                     
                     �    d                    
                    �    d                    
                    �    d                 
   
             
       �    d                    $
                    �    d                    $
                    �    d                    $
                    �    d                    *
                     �    e                     7
                     �    e                    A
                    �    e                    A
                    �    e                    A
                    �    e                    A
                    �    e                    A
                    �    e                    A
                    �    e                    A
                    �    e   %                 P
                     �    f                     ]
                     �    f   "                 s
                    �    f   (                 y
                     �    g                      z
                     5�_�                    h        ����                                                                                                                                                                                                                                                                                                                                                             f:w�     �   g   i   �       5��    g                      z
                     �    g                    �
                    5�_�                    h   #    ����                                                                                                                                                                                                                                                                                                                                                             f:w�     �   g   i   �      $            count => words_received,5��    g   #                  �
                     5�_�                    �        ����                                                                                                                                                                                                                                                                                                                                                             f:�     �   �   �   �                      encrypt_in�   �   �   �                      �   �   �   �    5��    �                      �                     �    �                      �                     �    �                      �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                 
   �             
       �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                 
   �             
       �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                 
   �             
       �    �          
          �      
              �    �                    �                    5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f:�&     �   �   �   �                      encrypt_in <= 5��    �                     �                     5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             f:�'     �   �   �   �                       encrypt_in <= ()5��    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    �    �                    �                    5�_�                    �   -    ����                                                                                                                                                                                                                                                                                                                                                             f:�)     �   �   �   �      -                encrypt_in <= (others => '0')5��    �   -                  �                     5�_�                    i   	    ����                                                                                                                                                                                                                                                                                                                                                             f:�?     �   i   l   �              �   i   k   �    5��    i                      �
              	       �    i                      �
                     �    i                     �
              	       �    j                      �
                     5�_�                    i       ����                                                                                                                                                                                                                                                                                                                                                             f:�E     �   h   j   �      
        );5��    h                     �
                     5�_�                    _       ����                                                                                                                                                                                                                                                                                                                                                             f:�I     �   ^   `   �      
        );5��    ^                     �	                     5�_�                    i       ����                                                                                                                                                                                                                                                                                                                                                             f:�K     �   i   l   �          �   i   k   �    5��    i                      �
                     �    i                      �
                     �    i                     �
                     �    j                     �
                     �    j                    �
                    �    j                     �
                     5�_�                    k       ����                                                                                                                                                                                                                                                                                                                                                             f:�b     �   k   m   �              port�   j   m   �          receiver_data: 5��    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                 
   �
             
       �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                    �
                    �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                    �
                    �    j                      �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                     �
                     �    j                    �
                    �    j                    �
                    �    j                    �
                    �    j   !                 �
                     �    k                     �
                     �    k                    �
                    �    k                    �
                    �    k                    �
                    5�_�                    l       ����                                                                                                                                                                                                                                                                                                                                                             f:�i     �   k   m   �              port map5��    k                     �
                     5�_�                    l       ����                                                                                                                                                                                                                                                                                                                                                             f:�n     �   k   m   �              port map()5��    k                     �
                     �    k                    �
                    �    k                    �
                    �    k                    �
                    �    k   &                 �
                    �    k   &                 �
                    �    k   &                 �
                    �    k   6                 �
                    �    k   6                 �
                    �    k   =                                     �    k   6                 �
                    �    k   6                 �
                    �    k   6                 �
                    �    k   E                  	                     5�_�                    l   E    ����                                                                                                                                                                                                                                                                                                                                                             f:�5     �   k   m   �      F        port map(reset, receiver_clk, done_receiving, received_data, )5��    k   E                  	                     �    k   F                 
                    5�_�                    l   M    ����                                                                                                                                                                                                                                                                                                                                                             f:�<     �   k   m   �      M        port map(reset, receiver_clk, done_receiving, received_data, message)5��    k   M                                       5�_�                     l   E    ����                                                                                                                                                                                                                                                                                                                                                             f:��     �   k   m   �      N        port map(reset, receiver_clk, done_receiving, received_data, message);5��    k   E                 	                    �    k   E              
   	             
       �    k   E       
          	      
              �    k   E              
   	             
       5�_�      !               q   N    ����                                                                                                                                                                                                                                                                                                                                                             f:��     �   p   q             encrypt_in <= received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data & received_data;5��    p                      3                    5�_�       "           !   p        ����                                                                                                                                                                                                                                                                                                                                                             f:��     �   o   p              -- received_data * 645��    o                                           5�_�   !   #           "   o        ����                                                                                                                                                                                                                                                                                                                                                             f:��     �   n   o           5��    n                                           5�_�   "   $           #   n        ����                                                                                                                                                                                                                                                                                                                                                             f:��     �   m   n           5��    m                                           5�_�   #   %           $   m        ����                                                                                                                                                                                                                                                                                                                                                             f:��     �   l   m           5��    l                                           5�_�   $   &           %   �        ����                                                                                                                                                                                                                                                                                                                                                             f:��     �   �   �          .                encrypt_in <= (others => '0');5��    �                      �      /               5�_�   %   (           &   �        ����                                                                                                                                                                                                                                                                                                                                                             f:��     �   �   �           5��    �                      �                     5�_�   &   )   '       (   �       ����                                                                                                                                                                                                                                                                                                                                                             f:�;     �   �   �   �      4                        if done_receiving = '1' then5��    �                    0                    �    �                     2                     �    �                     1                     �    �                    0                    �    �   -                  B                     �    �   ,                  A                     �    �   +                  @                     �    �   *                  ?                     �    �   )                  >                     �    �   (                  =                     �    �   '                  <                     �    �   &                  ;                     �    �   %                  :                     �    �   $                  9                     �    �   #                  8                     �    �   "                  7                     �    �   !                  6                     �    �                      5                     �    �                     4                     �    �                     3                     �    �                     2                     �    �                     1                     �    �                    0                    �    �                    0                    �    �                    0                    5�_�   (   *           )   C       ����                                                                                                                                                                                                                                                                                                                                                             f:��     �   C   E   �    �   C   D   �    5��    C                      W                      5�_�   )   +           *   D       ����                                                                                                                                                                                                                                                                                                                                                             f:��    �   C   E   �          signal done_receiving: bit;5��    C                     p                     �    C                     r                     �    C                     q                     �    C                     p                     �    C                     o                     �    C                     n                     �    C                     m                     �    C                     l                     �    C                     k                     �    C                     j                     �    C                     i                     �    C                     h                     �    C                     g                     �    C                     f                     �    C                     e                     �    C                     d                     �    C                     c                     �    C                    b                    �    C                    b                    �    C                    b                    5�_�   *   ,           +           ����                                                                                                                                                                                                                                                                                                                                                             f:��     �         �          end component�         �          component�         �          �         �    5��                          �                     �                          �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                     	   �             	       �              	          �      	              �                        �                    �                         �                     �                         �                     �                         �                     �                        �                    �                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �       #                  �                     �       "                  �                     �       !                  �                     �                          �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                         �                     �                        �                    �                        �                    �                        �                    �       $                 �                     �                         �                    �                         �                    �                                              �                                              �                                              �       
                                       �       	                                       �                     	                	       �              	                	              �                     
                
       5�_�   +   -           ,          ����                                                                                                                                                                                                                                                                                                                                                             f:��     �         �    �         �    5��                          �              �       5�_�   ,   .           -          ����                                                                                                                                                                                                                                                                                                                                                       f:��    �         �              MAX_COUNT: natural       );   
    port (   K        clk, rst, enable: in bit;                            -- Clock input           done: out bit;   B        count : out natural       -- 6-bit count output (64 steps)       );�         �          generic(5��                         �                     �                                              �                         .                     �                         9                     �                         H                     �                         �                     �                         �                     �                         �                     5�_�   -   /           .          ����                                                                                                                                                                                                                                                                                                                                                       f:��     �   !   #   �          end component�       #   �          component shift_reg_byte�      "   �          �      !   �    5��                                               �                                               �                                              �                                               �                         #                    �                         #                    �                         #                    �                         #                    �                         1                     �    !                     2                    �    !                     2                    �    !                     :                     �    !                 	   :             	       �    !          	          :      	              �    !                 
   :             
       5�_�   .   0           /   !       ����                                                                                                                                                                                                                                                                                                                                                       f:��     �   !   '   �    �   !   "   �    5��    !                      2              �       5�_�   /   1           0   "       ����                                                                                                                                                                                                                                                                                                                            "          &                 f:��    �   "   '   �      !        rst, clk, enable: in bit;   (        data: in bit_vector(7 downto 0);   '        q: out bit_vector(511 downto 0)       );�   !   #   �      
    port (5��    !                     6                     �    "                     E                     �    #                     k                     �    $                     �                     �    %                     �                     5�_�   0   2           1   V       ����                                                                                                                                                                                                                                                                                                                            "          &                 f:��     �   U   W   �          �   U   W   �    5��    U                      A                     �    U                  
   E              
       5�_�   1   3           2   V       ����                                                                                                                                                                                                                                                                                                                            "          &                 f:��     �   U   W   �          signal wor5��    U                     O                     5�_�   2   4           3   V       ����                                                                                                                                                                                                                                                                                                                            "          &                 f:��     �   U   X   �          signal wor[�   V   X              ]�   U   X   �          signal wor[]5��    U                    P                     �    U                    P                     �    V                      Q                     5�_�   3   5           4   W        ����                                                                                                                                                                                                                                                                                                                            "          &                 f:��     �   V   W                  ]5��    V                      Q                     5�_�   4   6           5   V       ����                                                                                                                                                                                                                                                                                                                            "          &                 f:��     �   U   W   �          signal wor[5��    U                    O                    �    U                    L                    �    U                    L                    �    U                    L                    5�_�   5   7           6   V       ����                                                                                                                                                                                                                                                                                                                            "          &                 f:��     �   U   W   �          signal words_received: nat5��    U                     _                     5�_�   6   8           7   V       ����                                                                                                                                                                                                                                                                                                                            "          &                 f:��    �   U   W   �           signal words_received: nat[]5��    U                    \                    �    U                    \                    �    U                    \                    5�_�   7   9           8   i       ����                                                                                                                                                                                                                                                                                                                            "          &                 f:�Z     �   h   j   �      $        port map(clock, sender_clk);5��    h                    �
                    �    h                    �
                    �    h                    �
                    �    h                    �
                    �    h                    �
                    �    h                    �
                    5�_�   8   :           9   h       ����                                                                                                                                                                                                                                                                                                                            "          &                 f:�p     �   g   i   �      K        generic map(5208) -- clock divido em 2 para judge e 5208 para placa5��    g                    ]
                    5�_�   9   ;           :   e       ����                                                                                                                                                                                                                                                                                                                            c          e          V       f:�t     �   b   f   �          receive_clk: slow_clk    K        generic map(1302)   -- Converte clock de 50M pra 19200Hz caso placa   &        port map(clock, receiver_clk);5��    b                     �	      �       �       5�_�   :   <           ;   b       ����                                                                                                                                                                                                                                                                                                                            c          e          V       f:�u    �   a   c   �      :    -- receiver_clk <= clock; -- Clock de 19200Hz do judge5��    a                     Z	      ;       8       5�_�   ;   =           <   h       ����                                                                                                                                                                                                                                                                                                                            c          e          V       f:�}    �   g   i   �      H        generic map(2) -- clock divido em 2 para judge e 5208 para placa5��    g          .           i
      .               5�_�   <   >           =   i       ����                                                                                                                                                                                                                                                                                                                            c          e          V       f:�    �   h   j   �      *        port map(receive_clk, sender_clk);5��    h                     �
                     5�_�   =   ?           >   h       ����                                                                                                                                                                                                                                                                                                                            c          e          V       f:�     �   g   i   �              generic map(2) -- 5��    g                    c
                    5�_�   >   @           ?   y       ����                                                                                                                                                                                                                                                                                                                            c          e          V       f:�k     �   x   z   �                   clk => receiver_clk,5��    x                    .                    �    x                    .                    �    x                    .                    �    x                    .                    5�_�   ?   A           @   y       ����                                                                                                                                                                                                                                                                                                                            c          e          V       f:�u   	 �   x   z   �                  clk => send_clk,5��    x                    .                    �    x                    .                    �    x                 
   .             
       �    x          
       
   .      
       
       �    x          
          .      
              �    x                 
   .             
       5�_�   @   B           A   �       ����                                                                                                                                                                                                                                                                                                                            c          e          V       f;[f   
 �   �   �   �      Q        port map(reset, receiver_clk, done_receiving, received_data, encrypt_in);5��    �                    	                    �    �                 
   	             
       �    �          
       
   	      
       
       �    �          
          	      
              �    �                 
   	             
       5�_�   A   C           B   �   2    ����                                                                                                                                                                                                                                                                                                                            c          e          V       f;`W     �   �   �   �      O        port map(reset, sender_clk, done_receiving, received_data, encrypt_in);5��    �   2                  #                     5�_�   B   D           C   �   7    ����                                                                                                                                                                                                                                                                                                                            c          e          V       f;``     �   �   �   �      T        port map(reset, sender_clk, done_receiving and , received_data, encrypt_in);5��    �   7                  (                     5�_�   C   E           D   �   8    ����                                                                                                                                                                                                                                                                                                                            c          e          V       f;`a     �   �   �   �      V        port map(reset, sender_clk, done_receiving and (), received_data, encrypt_in);5��    �   8                  )                     �    �   8                 )                    �    �   8                 )                    �    �   8                 )                    5�_�   D   F           E   �   @    ����                                                                                                                                                                                                                                                                                                                            c          e          V       f;`y    �   �   �   �      ^        port map(reset, sender_clk, done_receiving and (state = ), received_data, encrypt_in);5��    �   @                  1                     �    �   @              	   1             	       �    �   @       	          1      	              �    �   @              	   1             	       5�_�   E   G           F   W       ����                                                                                                                                                                                                                                                                                                                            c          e          V       f;`�     �   W   Y   �          �   W   Y   �    5��    W                      �                     �    W                     �                     �    W                    �                    5�_�   F   H           G   �       ����                                                                                                                                                                                                                                                                                                                            d          f          V       f;`�     �   �   �   �          �   �   �   �    5��    �                      �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    �    �                    �                    �    �                    �                    5�_�   G   I           H   �   $    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;`�     �   �   �   �      g        port map(reset, sender_clk, done_receiving and (state = receiving), received_data, encrypt_in);5��    �   $       &          J      &              �    �   $                 J                    �    �   $                 J                    �    �   $                 J                    5�_�   H   J           I   �       ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;`�     �   �   �   �          shift_message <= �   �   �   �    5��    �                  &                 &       5�_�   I   K           J   �   ;    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;`�    �   �   �   �      ;    shift_message <= done_receiving and (state = receiving)5��    �   ;                  )                     5�_�   J   L           K   �   $    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;`�    �   �   �   �      <    shift_message <= done_receiving and (state = receiving);5��    �   $                                     5�_�   K   M           L   �   $    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;a     �   �   �          :    shift_message <= done_receiving & (state = receiving);5��    �                      �      ;               5�_�   L   N           M   �        ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;a     �   �   �   �    �   �   �   �    5��    �                      f              ;       5�_�   M   O           N   �       ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;a     �   �   �   �      :    shift_message <= done_receiving & (state = receiving);5��    �                     j                     5�_�   N   P           O   �   !    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;a!     �   �   �   �      F                shift_message <= done_receiving & (state = receiving);5��    �   !       $           �      $               5�_�   O   Q           P   �   !    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;a"     �   �   �   �      "                shift_message <= ;5��    �   !                  �                     5�_�   P   S           Q   �   "    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;a#     �   �   �   �      $                shift_message <= '';5��    �   "                  �                     5�_�   Q   T   R       S   �   "    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;a0     �   �   �   �                                  �   �   �   �    5��    �                      <                     �    �                     X                     �    �                    X                    �    �                    X                    �    �                    X                    5�_�   S   U           T   �   -    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;a3     �   �   �   �      -                            shift_message <= 5��    �   -                  i                     5�_�   T   V           U   �   .    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;a4     �   �   �   �      /                            shift_message <= ''5��    �   .                  j                     5�_�   U   W           V   �   0    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;a5     �   �   �   �      0                            shift_message <= '1'5��    �   0                  l                     5�_�   V   X           W   �   /    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;aF     �   �   �   �                                  �   �   �   �    5��    �                      !                     �    �                     =                     �    �                    =                    �    �                    =                    �    �                    =                    5�_�   W   Y           X   �   -    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;aJ     �   �   �   �      -                            shift_message <= 5��    �   -                  N                     5�_�   X   Z           Y   �   .    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;aJ     �   �   �   �      /                            shift_message <= ''5��    �   .                  O                     5�_�   Y   [           Z   �   0    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;aK    �   �   �   �      0                            shift_message <= '0'5��    �   0                  Q                     5�_�   Z   \           [   �   .    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;a�    �   �   �   �      1                            shift_message <= '1';5��    �   -                 i                    �    �   -                 i                    �    �   -                 i                    �    �   -                 i                    �    �   -                 i                    �    �   -                 i                    �    �   -                 i                    �    �   -                 i                    5�_�   [   ]           \   �   %    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;bi     �   �   �          <                            shift_message <= done_receiving;5��    �                      <      =               5�_�   \   ^           ]   �        ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;bj     �   �   �   �    �   �   �   �    5��    �                      �              =       5�_�   ]   _           ^   �       ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;bl    �   �   �   �      <                            shift_message <= done_receiving;5��    �                     �                     5�_�   ^   `           _   x       ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;c6    �   w   y   �              generic map(64)5��    w                    %                    5�_�   _   a           `   �   #    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;g1     �   �   �   �      $            tx_done => done_sending,5��    �   #                  $                     5�_�   `   b           a   �        ����                                                                                                                                                                                                                                                                                                                            w   '                 V   '    f;g?     �   �   �   �    5��    �                      �              	       �    �                      �                     5�_�   a   c           b   �        ����                                                                                                                                                                                                                                                                                                                            w   '                 V   '    f;g?     �   �   �   �    �   �   �   �    5��    �               	       �              
      5�_�   b   d           c   �       ����                                                                                                                                                                                                                                                                                                                            �          �   	       v   	    f;gE     �   �   �   �      ,    receiver_counter: counter_generic_enable5��    �                    �                    5�_�   c   e           d   �       ����                                                                                                                                                                                                                                                                                                                            �          �   	       v   	    f;gM     �   �   �   �              generic map(65)5��    �                    �                    5�_�   d   f           e   �       ����                                                                                                                                                                                                                                                                                                                            �          �   	       v   	    f;gf     �   �   �   �      %            enable => done_receiving,5��    �          	          0      	              5�_�   e   g           f   �   #    ����                                                                                                                                                                                                                                                                                                                            �          �   	       v   	    f;gq     �   �   �   �      (            done => done_receiving_msgi,5��    �   #                 \                    5�_�   f   h           g   �       ����                                                                                                                                                                                                                                                                                                                            �          �   !       v   !    f;gy     �   �   �   �      (            done => done_receiving_haso,5��    �          	          R      	              5�_�   g   i           h   �   #    ����                                                                                                                                                                                                                                                                                                                            �          �   !       v   !    f;g     �   �   �   �      )            tx_done => done_sending_haso,5��    �   #                  $                     5�_�   h   j           i   �       ����                                                                                                                                                                                                                                                                                                                            �          �   !       v   !    f;g�     �   �   �   �      #            count => words_received5��    �                    v                    5�_�   i   k           j   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;i�     �   �   �   �    5��    �                      �                     �    �                      �                     5�_�   j   l           k   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;i�     �   �   �   �    �   �   �   �    5��    �                      �              q       5�_�   k   m           l   �       ����                                                                                                                                                                                                                                                                                                                            �          �          v       f;j      �   �   �   �      !    receiver_data: shift_reg_byte5��    �                    �                    5�_�   l   n           m   �       ����                                                                                                                                                                                                                                                                                                                            �          �          v       f;j     �   �   �   �          sender_data: shift_reg_byte5��    �                     �                     5�_�   m   o           n   �   $    ����                                                                                                                                                                                                                                                                                                                            �          �          v       f;j9     �   �   �   �      N        port map(reset, sender_clk, shift_message, received_data, encrypt_in);5��    �   $                 �                    5�_�   n   p           o   �   (    ����                                                                                                                                                                                                                                                                                                                            �          �          v       f;jG     �   �   �   �      I        port map(reset, sender_clk, get_data, received_data, encrypt_in);5��    �   (                  �                     �    �   ,                 �                    5�_�   o   q           p   �   8    ����                                                                                                                                                                                                                                                                                                                            �          �          v       f;jY     �   �   �   �      S        port map(reset, sender_clk, get_encrypted_data, received_data, encrypt_in);5��    �   8                 �                    �    �   8                 �                    �    �   8                 �                    �    �   8                 �                    5�_�   p   r           q   �   E    ����                                                                                                                                                                                                                                                                                                                            �          �          v       f;jh     �   �   �   �      Q        port map(reset, sender_clk, get_encrypted_data, encrypt_out, encrypt_in);5��    �   E       
          �      
              �    �   E                 �                    �    �   E                 �                    �    �   E                 �                    �    �   E                 �                    �    �   M                 �                    5�_�   q   s           r   �       ����                                                                                                                                                                                                                                                                                                                            �          �   *       v   *    f;ju    �   �   �   �      ,            data => encrypt_out(7 downto 0),5��    �                    :                    �    �                    :                    �    �                    :                    �    �                    :                    5�_�   r   t           s   W       ����                                                                                                                                                                                                                                                                                                                            �          �   *       v   *    f;j�     �   W   Y   �          �   W   Y   �    5��    W                      �                     �    W                     �                     �    W                    �                    �    W                    �                    �    W                    �                    �    W                    �                    �    W                    �                    �    W                    �                    �    W                    �                    5�_�   s   u           t   X       ����                                                                                                                                                                                                                                                                                                                            �          �   *       v   *    f;j�     �   Y   [   �      
    signal�   X   [   �          �   X   Z   �    5��    X                      �                     �    X                     �                     �    X                    �                    �    X                    �                    �    X                    �                    �    X                    �                    �    X                    �                    �    X                    �                    �    X   "                 �                     �    Y                     �                     �    Y                    �                    �    Y                    �                    �    Y                 
   �             
       �    Y                    �                    �    Y                 
   �             
       �    Y          
       
   �      
       
       �    Y          
          �      
              �    Y                    �                    �    Y                    �                    �    Y                    �                    �    Y                    �                    5�_�   t   v           u   '       ����                                                                                                                                                                                                                                                                                                                            �          �   *       v   *    f;j�     �   )   +   �          end component�   (   +   �          component�   '   *   �          �   '   )   �    5��    '                      �                     �    '                      �                     �    '                     �                     �    (                     �                     �    (                 	   �             	       �    (          	          �      	              �    (                    �                    �    (                    �                    �    (                    �                    �    (                    �                    �    (                     �                     �    )                                          �    )                                          �    )                                          �    )                 	                	       �    )          	                	              �    )                 
                
       5�_�   u   w           v   *       ����                                                                                                                                                                                                                                                                                                                            �          �   *       v   *    f;j�     �   )   /   �    �   *   +   �    5��    )                                     �       5�_�   v   x           w   *       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;j�    �   *   /   �      !        rst, clk, enable: in bit;   '        d: in bit_vector(255 downto 0);   %        q: out bit_vector(7 downto 0)       );�   )   +   �      
    port (5��    )                                          �    *                                          �    +                     9                     �    ,                     e                     �    -                     �                     5�_�   w   y           x   `       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k!     �   _   a   �          signal encrypt_byte: bit;5��    _                     l	                     �    _                 
   i	             
       �    _          
          i	      
              �    _                 
   i	             
       5�_�   x   z           y   `   #    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k#     �   _   a   �      $    signal encrypt_byte: bit_vector;5��    _   #                  s	                     5�_�   y   {           z   `   $    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k$     �   _   a   �      &    signal encrypt_byte: bit_vector();5��    _   $                  t	                     �    _   &                 v	                    �    _   &                 v	                    �    _   &                 v	                    5�_�   z   |           {   `       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k,     �   _   a   �      0    signal encrypt_byte: bit_vector(7 downto 0);5��    _                     b	                     5�_�   {   }           |   `       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k-     �   _   `          2    signal encrypted_byte: bit_vector(7 downto 0);5��    _                      P	      3               5�_�   |   ~           }   \        ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k.     �   [   ]   �    �   \   ]   �    5��    [                      �              3       5�_�   }              ~   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k5     �   �   �   �      !            data => encrypt_byte,5��    �                     �                     5�_�   ~   �              �   L    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k9    �   �   �   �      S        port map(reset, sender_clk, get_encrypted_data, encrypt_out, encrypt_byte);5��    �   L                  +                     5�_�      �           �   b       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;kO     �   b   d   �          �   b   d   �    5��    b                      �	                     �    b                  
   �	              
       �    b                    �	                    �    b                    �	                    �    b                    �	                    �    b                    �	                    5�_�   �   �           �   �   "    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;kb     �   �   �   �                                  �   �   �   �    5��    �                      G                     �    �                     c                     �    �                    c                    �    �                    c                    �    �                    c                    5�_�   �   �           �   �   0    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;ke     �   �   �   �      0                            get_encrypted_data <5��    �   0                  w                     5�_�   �   �           �   �   1    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;kf     �   �   �   �      2                            get_encrypted_data <''5��    �   0                 w                    5�_�   �   �           �   �   2    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;kg     �   �   �   �      2                            get_encrypted_data <= 5��    �   2                  y                     5�_�   �   �           �   �   3    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;kh     �   �   �   �      4                            get_encrypted_data <= ''5��    �   3                  z                     5�_�   �   �           �   �   5    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;ki     �   �   �   �      5                            get_encrypted_data <= '1'5��    �   5                  |                     5�_�   �   �           �   �   "    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;km     �   �   �   �                              �   �   �   �    5��    �                      �                     �    �                     �                    �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   �   .    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k�     �   �   �   �      .                        get_encrypted_data <= 5��    �   .                  �                     5�_�   �   �           �   �   /    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k�     �   �   �   �      0                        get_encrypted_data <= ''5��    �   /                  �                     5�_�   �   �           �   �   1    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k�     �   �   �   �      1                        get_encrypted_data <= '0'5��    �   1                  �                     5�_�   �   �           �   �   1    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k�     �   �   �          6                            get_encrypted_data <= '1';5��    �                      G      7               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k�     �   �   �   �    �   �   �   �    5��    �                      �              7       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k�     �   �   �   �      6                            get_encrypted_data <= '1';5��    �                     �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k�     �   �   �          2                        get_encrypted_data <= '0';5��    �                      �      3               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k�     �   �   �   �    �   �   �   �    5��    �                      z              3       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;k�    �   �   �   �      2                        get_encrypted_data <= '0';5��    �                     �                     5�_�   �   �           �   �   $    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;l     �   �   �          2                        get_encrypted_data <= '1';5��    �                      �      3               5�_�   �   �           �   �   $    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;l�     �   �   �   �    �   �   �   �    5��    �                      ~              3       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;l�     �   �   �   �      2                        get_encrypted_data <= '1';5��    �                     �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;l�     �   �   �          6                            get_encrypted_data <= '0';5��    �                      G      7               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;l�     �   �   �   �    �   �   �   �    5��    �                      �              7       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;l�    �   �   �   �      6                            get_encrypted_data <= '0';5��    �                     �                     5�_�   �   �           �   �   '    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;os     �   �   �          6                            get_encrypted_data <= '1';5��    �                      G      7               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;ow     �   �   �   �    �   �   �   �    5��    �                      �              7       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;ox    �   �   �   �      6                            get_encrypted_data <= '1';5��    �                     �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;o�     �   �   �          2                        get_encrypted_data <= '0';5��    �                      �      3               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;o�     �   �   �   �    �   �   �   �    5��    �                      z              3       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;o�    �   �   �   �      2                        get_encrypted_data <= '0';5��    �                     �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;p�     �   �   �   �                                  �   �   �   �    5��    �                      z                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   �   *    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;p�     �   �   �   �      *                            if rising_edge5��    �   *                  �                     5�_�   �   �           �   �   +    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;p�     �   �   �   �      ,                            if rising_edge()5��    �   +                  �                     �    �   +                 �                    �    �   +              
   �             
       �    �   +       
       
   �      
       
       �    �   +       
          �      
              �    �   +              
   �             
       5�_�   �   �           �   �   6    ����                                                                                                                                                                                                                                                                                                                            *          .                 f;p�     �   �   �   �      6                            if rising_edge(sender_clk)5��    �   6                  �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;p�     �   �   �   �      6                            get_encrypted_data <= '0';5��    �                     �                     5�_�   �   �   �       �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;p�    �   �   �   �                                       �   �   �   �    5��    �                      �              !       �    �                                           �    �                      �                     �    �                                           �    �   "                                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;qE    �   �   �   �          process(clock, reset) is5��    �                     k                     �    �                 
   m             
       �    �          
          m      
              �    �                 
   m             
       5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;q�     �   �   �          ;                            if rising_edge(sender_clk) then   :                                get_encrypted_data <= '0';   #                            end if;5��    �                      �      �               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;q�     �   �   �   �    �   �   �   �    5��    �                      �              �       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f;q�     �   �   �   �      ;                            if rising_edge(sender_clk) then5��    �                     �                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 f;q�     �   �   �   �      :                                get_encrypted_data <= '0';5��    �                                          5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 f;q�    �   �   �   �      #                            end if;5��    �                     R                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;r     �   �   �          7                        if rising_edge(sender_clk) then   6                            get_encrypted_data <= '0';                           end if;5��    �                      �      �               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;r     �   �   �   �    5��    �                      �                     �    �                     �                    �    �                      �                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;r     �   �   �   �    �   �   �   �    5��    �                      �              �       5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;r!     �   �   �           5��    �                      �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;r#     �   �   �   �      7                        if rising_edge(sender_clk) then5��    �                     �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;r%     �   �   �   �      6                            get_encrypted_data <= '0';5��    �                     �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;r&     �   �   �   �                              end if;5��    �                     �                     5�_�   �   �           �   �   #    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;r,    �   �   �   �      '        if rising_edge(sender_clk) then5��    �   #                  �                     �    �   '                 �                    �    �   (                 �                    �    �   (                 �                    �    �   (                 �                    �    �   (              	   �             	       �    �   0              	   �             	       5�_�   �   �           �   �   $    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;s&     �   �   �   �      U        port map(reset, sender_clk, get_encrypted_data, encrypt_out, encrypted_byte);5��    �   $                 '                    5�_�   �   �           �   �   "    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;sZ     �   �   �   �    �   �   �   �    5��    �                      E              9       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;s^     �   �   �   �      8                        shift_message <= done_receiving;5��    �                     c                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;s_     �   �   �   �      9                        shift__message <= done_receiving;5��    �                     c                     �    �                    ]                    �    �                    ]                    �    �                    ]                    5�_�   �   �           �   �   /    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;sb     �   �   �   �      J                        shift_encrypted_message_message <= done_receiving;5��    �   /       	           t      	               5�_�   �   �           �   �   /    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;sc     �   �   �   �      A                        shift_encrypted_message<= done_receiving;5��    �   /                  t                     5�_�   �   �           �   �   8    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;sg     �   �   �   �      B                        shift_encrypted_message <= done_receiving;5��    �   8       	          }      	              �    �   8                 }                    �    �   3       	          x      	              �    �   3                 x                    �    �   3                 x                    �    �   3                 x                    �    �   3                 x                    5�_�   �   �           �   �   $    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;s�     �   �   �   �                      �   �   �   �    5��    �                      �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   �   &    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;s�     �   �   �   �      &                aquire_sender_data <= 5��    �   &                                       5�_�   �   �           �   �   '    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;s�     �   �   �   �      (                aquire_sender_data <= ''5��    �   '                                       5�_�   �   �           �   �   )    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;s�     �   �   �   �      )                aquire_sender_data <= '0'5��    �   )                                       5�_�   �   �           �   �   )    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;s�     �   �   �   �    �   �   �   �    5��    �                      �              +       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;s�     �   �   �   �      *                aquire_sender_data <= '0';5��    �                     �                     5�_�   �   �           �   �   '    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;s�     �   �   �   �      N                        if done_sending then -- numero de stop bits arbitrario5��    �   '                  �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   �   +    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;s�     �   �   �   �                                  �   �   �   �    5��    �                      �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   �   7    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;t     �   �   �   �      7                            shift_encrypted_message <= 5��    �   7                                       5�_�   �   �           �   �   8    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;t     �   �   �   �      9                            shift_encrypted_message <= ''5��    �   8                                       5�_�   �   �           �   �   :    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;t     �   �   �   �      :                            shift_encrypted_message <= '0'5��    �   :                                       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;t     �   �   �   �      Z        port map(reset, sender_clk, shift_encrypted_message, encrypt_out, encrypted_byte);5��    �                                        �    �                                        �    �                                        �    �                                        5�_�   �   �           �   �   &    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;t5     �   �   �   �                              �   �   �   �    5��    �                      �                     �    �                     �                     �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   �   .    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;t:     �   �   �   �      .                        aquire_sender_data <= 5��    �   .                  �                     5�_�   �   �           �   �   /    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;t:     �   �   �   �      0                        aquire_sender_data <= ''5��    �   /                  �                     5�_�   �   �           �   �   1    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;t<     �   �   �   �      1                        aquire_sender_data <= '1'5��    �   1                  �                     �    �   2                  �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;tD     �   �   �   �      k        port map(not aquire_sender_data, sender_clk, shift_encrypted_message, encrypt_out, encrypted_byte);5��    �                                          5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;tT    �   �   �   �      &            get_encrypted_data <= '0';5��    �                    �                    �    �                    �                    �    �                    �                    �    �                    �                    5�_�   �   �           �   b       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;t�     �   c   e   �      
    signal�   b   e   �          �   b   d   �    5��    b                      �	                     �    b                  
   �	              
       �    b                    �	                    �    b                    �	                    �    b                    �	                    �    b   #                 �	                     �    c                     �	                     �    c                    �	                    �    c                    �	                    �    c                 
   �	             
       �    c                    �	                    �    c                    �	                    �    c                    �	                    5�_�   �   �           �   �   $    ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;t�     �   �   �   �    �   �   �   �    5��    �                      D              &       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;t�    �   �   �   �      %                shift_message <= '0';5��    �                    T                    �    �                    T                    �    �                    T                    �    �                    T                    5�_�   �   �           �   e       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;u     �   d   e          #    signal get_encrypted_data: bit;5��    d                      
      $               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;u    �   �   �          2                        get_encrypted_data <= '1';5��    �                      �      3               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;uZ     �   �   �          =        if rising_edge(sender_clk) and (state = sending) then5��    �                      �      >               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;u[     �   �   �                  end if;5��    �                      �                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;u\     �   �   �          &            aquire_sender_data <= '0';5��    �                      �      '               5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;u_     �   �   �   �    �   �   �   �    5��    �                      �              '       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       f;ua     �   �   �   �      &            aquire_sender_data <= '0';5��    �                     �                     5�_�   �   �           �   c        ����                                                                                                                                                                                                                                                                                                                                                             f;z�     �   c   e   �    �   c   d   �    5��    c                      �	              $       5�_�   �   �           �   d       ����                                                                                                                                                                                                                                                                                                                                                             f;z�     �   c   e   �      #    signal aquire_sender_data: bit;5��    c                    �	                    �    c                    �	                    �    c                    �	                    �    c                    �	                    �    c                    �	                    5�_�   �   �           �   d       ����                                                                                                                                                                                                                                                                                                                                                             f;z�     �   c   e   �      !    signal start_encrypting: bit;5��    c                     �	                     5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                                                             f;z�     �   �   �   �              �   �   �   �    5��    �                                           �    �                                           �    �                                        �    �                                        �    �                                          �    �                                          �    �                                          �    �                                        �    �                     +                     �    �                     *                     �    �                     )                     �    �                     (                     �    �                     '                     �    �                     &                     �    �                     %                     �    �                     $                     �    �                     #                     �    �                     "                     �    �                     !                     �    �                                           �    �                                          �    �   
                                       �    �   	                                       �    �                                          �    �                                          �    �                                          �    �                                          �    �                                        �    �                                        �    �                                        �    �   "                  6                     �    �   !                  5                     �    �                     4                    �    �                     4                    �    �                     4                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                             f;z�     �   �   �   �      (            rst => not start_encrypting,5��    �                    �                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             f;{     �          �    �         �    5��                                           (       5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             f;{   ! �         �    5��                          (                      5�_�   �   �           �   �   ,    ����                                                                                                                                                                                                                                                                                                                                                             f;{%     �   �   �   �      S                        if done_sending_haso then -- numero de stop bits arbitrario5��    �   ,                  �                     5�_�   �   �           �   �   -    ����                                                                                                                                                                                                                                                                                                                                                             f;{%     �   �   �   �      T                        if done_sending_haso  then -- numero de stop bits arbitrario5��    �   -                  �                     5�_�   �   �           �   �   .    ����                                                                                                                                                                                                                                                                                                                                                             f;{&     �   �   �   �      V                        if done_sending_haso '' then -- numero de stop bits arbitrario5��    �   -                  �                     �    �   -                 �                    5�_�   �   �           �   �   /    ����                                                                                                                                                                                                                                                                                                                                                             f;{'     �   �   �   �      V                        if done_sending_haso =  then -- numero de stop bits arbitrario5��    �   /                  �                     5�_�   �   �           �   �   0    ����                                                                                                                                                                                                                                                                                                                                                             f;{(   " �   �   �   �      X                        if done_sending_haso = '' then -- numero de stop bits arbitrario5��    �   0                  �                     5�_�   �   �           �   t        ����                                                                                                                                                                                                                                                                                                                                                  V        f=&v     �   s   u   �      7    receiver_clk <= clock; -- Clock de 19200Hz do judge5��    s                     V      8       ;       5�_�   �   �           �   w        ����                                                                                                                                                                                                                                                                                                                            u           w           V        f=&x   # �   t   x   �          -- receive_clk: slow_clk    N    --     generic map(1302)   -- Converte clock de 50M pra 19200Hz caso placa   )    --     port map(clock, receiver_clk);5��    t                     �      �       �       5�_�   �   �           �   w        ����                                                                                                                                                                                                                                                                                                                            u           w           V        fB��     �   t   x   �          receive_clk: slow_clk    K        generic map(1302)   -- Converte clock de 50M pra 19200Hz caso placa   &        port map(clock, receiver_clk);5��    t                     �      �       �       5�_�   �   �           �   t        ����                                                                                                                                                                                                                                                                                                                            u           w           V        fB��   $ �   s   u   �      :    -- receiver_clk <= clock; -- Clock de 19200Hz do judge5��    s                     V      ;       8       5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB��     �   �   �   �                              �   �   �   �    5��    �                      �                     �    �                      �                     �    �                     �                     �    �                    �                    5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB��     �   �   �                                  when 5��    �                      �                     5�_�   �   �   �       �   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB�[     �   �   �   �      (    process(clock, sender_clk, reset) is5��    �                     "                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB�[     �   �   �   �      #    process(, sender_clk, reset) is5��    �                     "                     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB�]   & �   �   �   �      "        if rising_edge(clock) then5��    �                    Y                    �    �                     `                     �    �                     _                     �    �                     ^                     �    �                     ]                     �    �                     \                     �    �                     [                     �    �                     Z                     �    �                 
   Y             
       �    �          
          Y      
              �    �                 
   Y             
       5�_�   �   �           �   t        ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB��     �   s   u   �      7    receiver_clk <= clock; -- Clock de 19200Hz do judge5��    s                     V      8       ;       5�_�   �   �           �   w        ����                                                                                                                                                                                                                                                                                                                            u          w           V        fB��   ' �   t   x   �          -- receive_clk: slow_clk    N    --     generic map(1302)   -- Converte clock de 50M pra 19200Hz caso placa   )    --     port map(clock, receiver_clk);5��    t                     �      �       �       5�_�   �   �           �   w        ����                                                                                                                                                                                                                                                                                                                            u          w           V        fC^Q     �   t   x   �          receive_clk: slow_clk    K        generic map(1302)   -- Converte clock de 50M pra 19200Hz caso placa   &        port map(clock, receiver_clk);5��    t                     �      �       �       5�_�   �   �           �   t        ����                                                                                                                                                                                                                                                                                                                            u          w           V        fC^S   ( �   s   u   �      :    -- receiver_clk <= clock; -- Clock de 19200Hz do judge5��    s                     V      ;       8       5�_�   �   �           �   t       ����                                                                                                                                                                                                                                                                                                                            u          w           V        fC`�     �   s   u   �      7    receiver_clk <= clock; -- Clock de 19200Hz do judge5��    s                     V      8       ;       5�_�   �   �           �   w       ����                                                                                                                                                                                                                                                                                                                            u          w          V       fC`�     �   t   x   �          -- receive_clk: slow_clk    N    --     generic map(1302)   -- Converte clock de 50M pra 19200Hz caso placa   )    --     port map(clock, receiver_clk);5��    t                     �      �       �       5�_�   �   �           �   v   9    ����                                                                                                                                                                                                                                                                                                                            v   9       v   ;       v   ;    fC`�     �   u   w   �      K        generic map(1302)   -- Converte clock de 50M pra 19200Hz caso placa5��    u   9                 �                    5�_�   �   �           �   v   ;    ����                                                                                                                                                                                                                                                                                                                            v   9       v   ;       v   ;    fC`�     �   u   w   �      K        generic map(1302)   -- Converte clock de 50M pra 20000Hz caso placa5��    u   ;                 �                    5�_�   �   �           �   v       ����                                                                                                                                                                                                                                                                                                                            v   9       v   ;       v   ;    fC`�   ) �   u   w   �      I        generic map(1302)   -- Converte clock de 50M pra 20kHz caso placa5��    u                    �                    5�_�   �   �           �   w       ����                                                                                                                                                                                                                                                                                                                            u          w          V       fCa�     �   t   x   �          receive_clk: slow_clk    I        generic map(1250)   -- Converte clock de 50M pra 20kHz caso placa   &        port map(clock, receiver_clk);5��    t                     �      �       �       5�_�   �              �   t       ����                                                                                                                                                                                                                                                                                                                            u          w          V       fCa�   * �   s   u   �      :    -- receiver_clk <= clock; -- Clock de 19200Hz do judge5��    s                     V      ;       8       5�_�   �                t       ����                                                                                                                                                                                                                                                                                                                            u          w          V       fCb�     �   s   u   �      7    receiver_clk <= clock; -- Clock de 19200Hz do judge5��    s                     V      8       ;       5�_�                  w       ����                                                                                                                                                                                                                                                                                                                            u          w          V       fCb�   + �   t   x   �          -- receive_clk: slow_clk    L    --     generic map(1250)   -- Converte clock de 50M pra 20kHz caso placa   )    --     port map(clock, receiver_clk);5��    t                     �      �       �       5�_�                 v       ����                                                                                                                                                                                                                                                                                                                            u          w          V       fCl	   , �   u   w   �      I        generic map(1250)   -- Converte clock de 50M pra 20kHz caso placa5��    u                    �                    5�_�                 v       ����                                                                                                                                                                                                                                                                                                                            u          w          V       fC�A     �   u   w   �      I        generic map(1249)   -- Converte clock de 50M pra 20kHz caso placa5��    u                    �                    5�_�                 v   I    ����                                                                                                                                                                                                                                                                                                                            u          w          V       fC�C     �   u   w   �      I        generic map(1250)   -- Converte clock de 50M pra 20kHz caso placa5��    u   I               "   �              "       5�_�                 v   k    ����                                                                                                                                                                                                                                                                                                                            u          w          V       fC�P   - �   u   w   �      k        generic map(1250)   -- Converte clock de 50M pra 20kHz caso placa, erro proposital de 1250 e n 12495��    u   k                                       5�_�                 l       ����                                                                                                                                                                                                                                                                                                                            u          w          V       fC��     �   l   n   �    �   l   m   �    5��    l                      �
                     5�_�                 m       ����                                                                                                                                                                                                                                                                                                                            v          x          V       fC��     �   l   n   �          signal done_sending: bit;5��    l                    �
                    5�_�                   �       ����                                                                                                                                                                                                                                                                                                                            v          x          V       fC��   . �   �   �   �                  reset => reset,5��    �                    e                    �    �                     h                     �    �                     g                     �    �                     f                     �    �                    e                    �    �                    e                    �    �                    e                    5�_�   �   �       �   �   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB�F     �   �   �   �                              �   �   �   �          ,                    when buffering_signal =>   &                        if rising_edge�   �   �   �      &                        if rising_edge5��    �                      �                     �    �                      �                     �    �                     �                     �    �                    �                    �    �                     �                     �    �                    �                    �    �                      �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                     �                     �    �                    �                    �    �   ,                 �                     �    �                     �                    �    �                                          �    �                                          �    �                                        �    �                                        �    �                                        5�_�   �   �           �   �   &    ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB�b     �   �   �   �      (                        if rising_edge()5��    �   &                                       5�_�   �   �           �   �   '    ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB�c     �   �   �   �      2                        if rising_edge(sender_clk)5��    �   '                                       �    �   '                                     �    �   '                                     �    �   '                                     �    �   *                                     �    �   '              
                
       �    �   '       
                
              �    �   '              
                
       5�_�   �   �           �   �   2    ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB�k     �   �   �   �      7                        if rising_edge(sender_clk) then   !                            state�   �   �   �      -                            state <= sending;   .                            aquire_sender_data�   �   �   �      2                            aquire_sender_data <= 5��    �   2                                       �    �   6                  !                     �    �   5                                        �    �   4                                       �    �   3                                     �    �   3                                     �    �   3                                     �    �   7                 "                     �    �                     #                    �    �                    A                    �    �                     A                     �    �                     @                     �    �                    ?                    �    �                    ?                    �    �                    ?                    �    �   %                 H                    �    �   %                 H                    �    �   %                 H                    �    �   -                 P                     �    �                     m                     �    �                     o                     �    �                     n                     �    �                    m                    �    �                    m                    �    �                    m                    5�_�   �   �           �   �   2    ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB�     �   �   �   �      4                            aquire_sender_data <= ''5��    �   2                  �                     5�_�   �   �           �   �   3    ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB��     �   �   �   �      5                            aquire_sender_data <= '0'5��    �   3                  �                     5�_�   �   �           �   �   5    ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB��     �   �   �   �      6                            aquire_sender_data <= '0';5��    �   5                  �                     5�_�   �   �           �   �   6    ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB��     �   �   �   �      6                            aquire_sender_data <= '0';                           end if;5��    �   6                 �                     �    �                    �                    �    �                    �                    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB��     �   �   �        5��    �                            3               5�_�   �   �           �   �   %    ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB��     �   �   �   �      6                            state <= buffering_signal;5��    �   %                 a                    �    �   (                  d                     �    �   '                  c                     �    �   &                  b                     �    �   %                 a                    �    �   %                 a                    �    �   %                 a                    5�_�   �               �   W   6    ����                                                                                                                                                                                                                                                                                                                            �           �           V        fB��   % �   V   X   �      O    type sha_state is (receiving, sending, encrypting, buffering_signal, idle);5��    V   6                  
                     �    V   7                                       �    V   6                 
                    �    V   7                                     �    V   7                                     �    V   7                                     5�_�   �           �   �   �       ����                                                                                                                                                                                                                                                                                                                            *          .                 f;p�     �   �   �   �    �   �   �   �      2                        get_encrypted_data <= '0';5��    �                      �              3       5�_�   Q           S   R   �   "    ����                                                                                                                                                                                                                                                                                                                            �   $       �   I       v   I    f;a,     �   �   �   �       5��    �                      <                     �    �                      <                     5�_�   &           (   '   �       ����                                                                                                                                                                                                                                                                                                                                                             f:�/     �   �   �   �      9                        if done_receiving_msgi = '1' then5��    �                                        �    �                                           �    �                                          �    �                                          �    �                                          �    �                                          �    �                                        �    �                                        �    �                                        5��