Vim�UnDo� %�d�+�:?�?D�4��c�Ϛp���^Ag   B                                   e��#    _�                             ����                                                                                                                                                                                                                                                                                                                                                             e��!     �                   �               5��                   B                      �      5�_�                             ����                                                                                                                                                                                                                                                                                                                                                             e��"    �                  5��                                                  5��