Vim�UnDo� o�����%��=O�g��D�<���~�z�%Q�1�n   �                                   f)$�    _�                     6        ����                                                                                                                                                                                                                                                                                                                                                             f(<�     �   5   6          		  par: out bit;5��    5                      �                     5�_�                    j       ����                                                                                                                                                                                                                                                                                                                                                             f(<�     �   i   j          					 par <= '0';5��    i                      �
                     5�_�                    �   
    ����                                                                                                                                                                                                                                                                                                                                                             f(<�     �   �   �          *									 par <= not data_to_parity(word);5��    �                      �      +               5�_�                            ����                                                                                                                                                                                                                                                                                                                                      '           V       f(<�    �              '   library IEEE;   use IEEE.NUMERIC_BIT.ALL;       entity counter_generic is       generic(           MAX_COUNT: natural       );   
    port (   J        clk, rst, start: in bit;                            -- Clock input           done: out bit;   B        count : out natural       -- 6-bit count output (64 steps)       );   end counter_generic;       -architecture Behavioral of counter_generic is   !    signal counter: natural := 0;       begin          &    counting: process(clk, rst, start)   	    begin           if rst = '1' then               counter <= 0;               done <= '0';   #        elsif rising_edge(clk) then   )            if counter = MAX_COUNT-1 then                   done <= '1';                   counter <= 0;               end if;   \            if (counter > 0 and counter < MAX_COUNT-1) or (start = '1' and counter = 0) then   '                counter <= counter + 1;               end if;           end if;       end process counting;           count <= counter;          end architecture;    5��            '                       �              5�_�                       0    ����                                                                                                                                                                                                                                                                                                                                                             f(m    �         �      0        data : in bit_vector(WIDTH-1 downto 0);5��       /                  M                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f(�A     �         �      entity serial_out is5��              
          0       
              5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f(�F     �         �      end serial_out;5��              
          p      
              5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                             f(�J     �         �      end sender;5��                        p                    5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                             f(�M     �         �      (architecture Behavioral of serial_out is5��              
          �      
              5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                             f(�R     �                        PARITY : natural := 1;5��                          �                      5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                             f(�S    �                #        POLARITY : boolean := TRUE;5��                          G       $               5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             f(��     �         �      M    function data_to_parity(data: bit_vector(WIDTH-1 downto 0)) return bit is5��                         �                     5�_�                       $    ����                                                                                                                                                                                                                                                                                                                                                             f(��     �          �      ,        variable xor_result: bit := data(0);5��       $                  
                     5�_�                    "   )    ����                                                                                                                                                                                                                                                                                                                                                             f(��    �   !   #   �      1            xor_result := xor_result xor data(i);5��    !   )                  j                     5�_�                    ?       ����                                                                                                                                                                                                                                                                                                                                                             f(��     �   >   @   �                      tx_done <= '1';5��    >                    �                    5�_�                    @   !    ����                                                                                                                                                                                                                                                                                                                                                             f(��     �   ?   A   �      !                serial_o <= '1';5��    ?                                           5�_�                    L   $    ����                                                                                                                                                                                                                                                                                                                                                             f(��     �   K   L          +                            tx_done <= '0';5��    K                      ?      ,               5�_�                    J   $    ����                                                                                                                                                                                                                                                                                                                                                             f(��     �   I   K   �    �   J   K   �    5��    I                      �              ,       5�_�                    J       ����                                                                                                                                                                                                                                                                                                                                                             f(��     �   I   K   �      +                            tx_done <= '0';5��    I                     �                     5�_�                    J       ����                                                                                                                                                                                                                                                                                                                                                             f(��     �   J   L   �    5��    J                                           �    J                                           5�_�                    y   #    ����                                                                                                                                                                                                                                                                                                                                                             f(�    �   y   {   �    �   y   z   �    5��    y                      t              0       5�_�                    j        ����                                                                                                                                                                                                                                                                                                                                                             f)$�     �   i   j          /                                tx_done <= '1';5��    i                      �      0               5�_�                    m       ����                                                                                                                                                                                                                                                                                                                                                             f)$�     �   m   o   �    �   m   n   �    5��    m                      p              0       5�_�                    n        ����                                                                                                                                                                                                                                                                                                                                                             f)$�     �   m   o   �      /                                tx_done <= '1';5��    m                     �                     5�_�                     i       ����                                                                                                                                                                                                                                                                                                                                                             f)$�    �   h   i          B                            if stop_bits_sent = (STOP_BITS-1) then   #                            end if;5��    h                      �      g               5��